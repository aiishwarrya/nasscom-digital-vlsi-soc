module picorv32a (clk,
    resetn,
    trap,
    mem_valid,
    mem_instr,
    mem_ready,
    mem_addr,
    mem_wdata,
    mem_wstrb,
    mem_rdata,
    mem_la_read,
    mem_la_write,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    pcpi_valid,
    pcpi_insn,
    pcpi_rs1,
    pcpi_rs2,
    pcpi_wr,
    pcpi_rd,
    pcpi_wait,
    pcpi_ready,
    irq,
    eoi,
    trace_valid,
    trace_data);
 input clk;
 input resetn;
 output trap;
 output mem_valid;
 output mem_instr;
 input mem_ready;
 output [31:0] mem_addr;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;
 input [31:0] mem_rdata;
 output mem_la_read;
 output mem_la_write;
 output [31:0] mem_la_addr;
 output [31:0] mem_la_wdata;
 output [3:0] mem_la_wstrb;
 output pcpi_valid;
 output [31:0] pcpi_insn;
 output [31:0] pcpi_rs1;
 output [31:0] pcpi_rs2;
 input pcpi_wr;
 input [31:0] pcpi_rd;
 input pcpi_wait;
 input pcpi_ready;
 input [31:0] irq;
 output [31:0] eoi;
 output trace_valid;
 output [35:0] trace_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire \alu_add_sub[0] ;
 wire \alu_add_sub[10] ;
 wire \alu_add_sub[11] ;
 wire \alu_add_sub[12] ;
 wire \alu_add_sub[13] ;
 wire \alu_add_sub[14] ;
 wire \alu_add_sub[15] ;
 wire \alu_add_sub[16] ;
 wire \alu_add_sub[17] ;
 wire \alu_add_sub[18] ;
 wire \alu_add_sub[19] ;
 wire \alu_add_sub[1] ;
 wire \alu_add_sub[20] ;
 wire \alu_add_sub[21] ;
 wire \alu_add_sub[22] ;
 wire \alu_add_sub[23] ;
 wire \alu_add_sub[24] ;
 wire \alu_add_sub[25] ;
 wire \alu_add_sub[26] ;
 wire \alu_add_sub[27] ;
 wire \alu_add_sub[28] ;
 wire \alu_add_sub[29] ;
 wire \alu_add_sub[2] ;
 wire \alu_add_sub[30] ;
 wire \alu_add_sub[31] ;
 wire \alu_add_sub[3] ;
 wire \alu_add_sub[4] ;
 wire \alu_add_sub[5] ;
 wire \alu_add_sub[6] ;
 wire \alu_add_sub[7] ;
 wire \alu_add_sub[8] ;
 wire \alu_add_sub[9] ;
 wire alu_eq;
 wire alu_lts;
 wire alu_ltu;
 wire \alu_out[0] ;
 wire \alu_out[10] ;
 wire \alu_out[11] ;
 wire \alu_out[12] ;
 wire \alu_out[13] ;
 wire \alu_out[14] ;
 wire \alu_out[15] ;
 wire \alu_out[16] ;
 wire \alu_out[17] ;
 wire \alu_out[18] ;
 wire \alu_out[19] ;
 wire \alu_out[1] ;
 wire \alu_out[20] ;
 wire \alu_out[21] ;
 wire \alu_out[22] ;
 wire \alu_out[23] ;
 wire \alu_out[24] ;
 wire \alu_out[25] ;
 wire \alu_out[26] ;
 wire \alu_out[27] ;
 wire \alu_out[28] ;
 wire \alu_out[29] ;
 wire \alu_out[2] ;
 wire \alu_out[30] ;
 wire \alu_out[31] ;
 wire \alu_out[3] ;
 wire \alu_out[4] ;
 wire \alu_out[5] ;
 wire \alu_out[6] ;
 wire \alu_out[7] ;
 wire \alu_out[8] ;
 wire \alu_out[9] ;
 wire \alu_out_q[0] ;
 wire \alu_out_q[10] ;
 wire \alu_out_q[11] ;
 wire \alu_out_q[12] ;
 wire \alu_out_q[13] ;
 wire \alu_out_q[14] ;
 wire \alu_out_q[15] ;
 wire \alu_out_q[16] ;
 wire \alu_out_q[17] ;
 wire \alu_out_q[18] ;
 wire \alu_out_q[19] ;
 wire \alu_out_q[1] ;
 wire \alu_out_q[20] ;
 wire \alu_out_q[21] ;
 wire \alu_out_q[22] ;
 wire \alu_out_q[23] ;
 wire \alu_out_q[24] ;
 wire \alu_out_q[25] ;
 wire \alu_out_q[26] ;
 wire \alu_out_q[27] ;
 wire \alu_out_q[28] ;
 wire \alu_out_q[29] ;
 wire \alu_out_q[2] ;
 wire \alu_out_q[30] ;
 wire \alu_out_q[31] ;
 wire \alu_out_q[3] ;
 wire \alu_out_q[4] ;
 wire \alu_out_q[5] ;
 wire \alu_out_q[6] ;
 wire \alu_out_q[7] ;
 wire \alu_out_q[8] ;
 wire \alu_out_q[9] ;
 wire \alu_shl[0] ;
 wire \alu_shl[10] ;
 wire \alu_shl[11] ;
 wire \alu_shl[12] ;
 wire \alu_shl[13] ;
 wire \alu_shl[14] ;
 wire \alu_shl[15] ;
 wire \alu_shl[16] ;
 wire \alu_shl[17] ;
 wire \alu_shl[18] ;
 wire \alu_shl[19] ;
 wire \alu_shl[1] ;
 wire \alu_shl[20] ;
 wire \alu_shl[21] ;
 wire \alu_shl[22] ;
 wire \alu_shl[23] ;
 wire \alu_shl[24] ;
 wire \alu_shl[25] ;
 wire \alu_shl[26] ;
 wire \alu_shl[27] ;
 wire \alu_shl[28] ;
 wire \alu_shl[29] ;
 wire \alu_shl[2] ;
 wire \alu_shl[30] ;
 wire \alu_shl[31] ;
 wire \alu_shl[3] ;
 wire \alu_shl[4] ;
 wire \alu_shl[5] ;
 wire \alu_shl[6] ;
 wire \alu_shl[7] ;
 wire \alu_shl[8] ;
 wire \alu_shl[9] ;
 wire \alu_shr[0] ;
 wire \alu_shr[10] ;
 wire \alu_shr[11] ;
 wire \alu_shr[12] ;
 wire \alu_shr[13] ;
 wire \alu_shr[14] ;
 wire \alu_shr[15] ;
 wire \alu_shr[16] ;
 wire \alu_shr[17] ;
 wire \alu_shr[18] ;
 wire \alu_shr[19] ;
 wire \alu_shr[1] ;
 wire \alu_shr[20] ;
 wire \alu_shr[21] ;
 wire \alu_shr[22] ;
 wire \alu_shr[23] ;
 wire \alu_shr[24] ;
 wire \alu_shr[25] ;
 wire \alu_shr[26] ;
 wire \alu_shr[27] ;
 wire \alu_shr[28] ;
 wire \alu_shr[29] ;
 wire \alu_shr[2] ;
 wire \alu_shr[30] ;
 wire \alu_shr[31] ;
 wire \alu_shr[3] ;
 wire \alu_shr[4] ;
 wire \alu_shr[5] ;
 wire \alu_shr[6] ;
 wire \alu_shr[7] ;
 wire \alu_shr[8] ;
 wire \alu_shr[9] ;
 wire alu_wait;
 wire \count_cycle[0] ;
 wire \count_cycle[10] ;
 wire \count_cycle[11] ;
 wire \count_cycle[12] ;
 wire \count_cycle[13] ;
 wire \count_cycle[14] ;
 wire \count_cycle[15] ;
 wire \count_cycle[16] ;
 wire \count_cycle[17] ;
 wire \count_cycle[18] ;
 wire \count_cycle[19] ;
 wire \count_cycle[1] ;
 wire \count_cycle[20] ;
 wire \count_cycle[21] ;
 wire \count_cycle[22] ;
 wire \count_cycle[23] ;
 wire \count_cycle[24] ;
 wire \count_cycle[25] ;
 wire \count_cycle[26] ;
 wire \count_cycle[27] ;
 wire \count_cycle[28] ;
 wire \count_cycle[29] ;
 wire \count_cycle[2] ;
 wire \count_cycle[30] ;
 wire \count_cycle[31] ;
 wire \count_cycle[32] ;
 wire \count_cycle[33] ;
 wire \count_cycle[34] ;
 wire \count_cycle[35] ;
 wire \count_cycle[36] ;
 wire \count_cycle[37] ;
 wire \count_cycle[38] ;
 wire \count_cycle[39] ;
 wire \count_cycle[3] ;
 wire \count_cycle[40] ;
 wire \count_cycle[41] ;
 wire \count_cycle[42] ;
 wire \count_cycle[43] ;
 wire \count_cycle[44] ;
 wire \count_cycle[45] ;
 wire \count_cycle[46] ;
 wire \count_cycle[47] ;
 wire \count_cycle[48] ;
 wire \count_cycle[49] ;
 wire \count_cycle[4] ;
 wire \count_cycle[50] ;
 wire \count_cycle[51] ;
 wire \count_cycle[52] ;
 wire \count_cycle[53] ;
 wire \count_cycle[54] ;
 wire \count_cycle[55] ;
 wire \count_cycle[56] ;
 wire \count_cycle[57] ;
 wire \count_cycle[58] ;
 wire \count_cycle[59] ;
 wire \count_cycle[5] ;
 wire \count_cycle[60] ;
 wire \count_cycle[61] ;
 wire \count_cycle[62] ;
 wire \count_cycle[63] ;
 wire \count_cycle[6] ;
 wire \count_cycle[7] ;
 wire \count_cycle[8] ;
 wire \count_cycle[9] ;
 wire \count_instr[0] ;
 wire \count_instr[10] ;
 wire \count_instr[11] ;
 wire \count_instr[12] ;
 wire \count_instr[13] ;
 wire \count_instr[14] ;
 wire \count_instr[15] ;
 wire \count_instr[16] ;
 wire \count_instr[17] ;
 wire \count_instr[18] ;
 wire \count_instr[19] ;
 wire \count_instr[1] ;
 wire \count_instr[20] ;
 wire \count_instr[21] ;
 wire \count_instr[22] ;
 wire \count_instr[23] ;
 wire \count_instr[24] ;
 wire \count_instr[25] ;
 wire \count_instr[26] ;
 wire \count_instr[27] ;
 wire \count_instr[28] ;
 wire \count_instr[29] ;
 wire \count_instr[2] ;
 wire \count_instr[30] ;
 wire \count_instr[31] ;
 wire \count_instr[32] ;
 wire \count_instr[33] ;
 wire \count_instr[34] ;
 wire \count_instr[35] ;
 wire \count_instr[36] ;
 wire \count_instr[37] ;
 wire \count_instr[38] ;
 wire \count_instr[39] ;
 wire \count_instr[3] ;
 wire \count_instr[40] ;
 wire \count_instr[41] ;
 wire \count_instr[42] ;
 wire \count_instr[43] ;
 wire \count_instr[44] ;
 wire \count_instr[45] ;
 wire \count_instr[46] ;
 wire \count_instr[47] ;
 wire \count_instr[48] ;
 wire \count_instr[49] ;
 wire \count_instr[4] ;
 wire \count_instr[50] ;
 wire \count_instr[51] ;
 wire \count_instr[52] ;
 wire \count_instr[53] ;
 wire \count_instr[54] ;
 wire \count_instr[55] ;
 wire \count_instr[56] ;
 wire \count_instr[57] ;
 wire \count_instr[58] ;
 wire \count_instr[59] ;
 wire \count_instr[5] ;
 wire \count_instr[60] ;
 wire \count_instr[61] ;
 wire \count_instr[62] ;
 wire \count_instr[63] ;
 wire \count_instr[6] ;
 wire \count_instr[7] ;
 wire \count_instr[8] ;
 wire \count_instr[9] ;
 wire \cpu_state[0] ;
 wire \cpu_state[1] ;
 wire \cpu_state[2] ;
 wire \cpu_state[3] ;
 wire \cpu_state[4] ;
 wire \cpu_state[5] ;
 wire \cpu_state[6] ;
 wire \cpuregs[0][0] ;
 wire \cpuregs[0][10] ;
 wire \cpuregs[0][11] ;
 wire \cpuregs[0][12] ;
 wire \cpuregs[0][13] ;
 wire \cpuregs[0][14] ;
 wire \cpuregs[0][15] ;
 wire \cpuregs[0][16] ;
 wire \cpuregs[0][17] ;
 wire \cpuregs[0][18] ;
 wire \cpuregs[0][19] ;
 wire \cpuregs[0][1] ;
 wire \cpuregs[0][20] ;
 wire \cpuregs[0][21] ;
 wire \cpuregs[0][22] ;
 wire \cpuregs[0][23] ;
 wire \cpuregs[0][24] ;
 wire \cpuregs[0][25] ;
 wire \cpuregs[0][26] ;
 wire \cpuregs[0][27] ;
 wire \cpuregs[0][28] ;
 wire \cpuregs[0][29] ;
 wire \cpuregs[0][2] ;
 wire \cpuregs[0][30] ;
 wire \cpuregs[0][31] ;
 wire \cpuregs[0][3] ;
 wire \cpuregs[0][4] ;
 wire \cpuregs[0][5] ;
 wire \cpuregs[0][6] ;
 wire \cpuregs[0][7] ;
 wire \cpuregs[0][8] ;
 wire \cpuregs[0][9] ;
 wire \cpuregs[10][0] ;
 wire \cpuregs[10][10] ;
 wire \cpuregs[10][11] ;
 wire \cpuregs[10][12] ;
 wire \cpuregs[10][13] ;
 wire \cpuregs[10][14] ;
 wire \cpuregs[10][15] ;
 wire \cpuregs[10][16] ;
 wire \cpuregs[10][17] ;
 wire \cpuregs[10][18] ;
 wire \cpuregs[10][19] ;
 wire \cpuregs[10][1] ;
 wire \cpuregs[10][20] ;
 wire \cpuregs[10][21] ;
 wire \cpuregs[10][22] ;
 wire \cpuregs[10][23] ;
 wire \cpuregs[10][24] ;
 wire \cpuregs[10][25] ;
 wire \cpuregs[10][26] ;
 wire \cpuregs[10][27] ;
 wire \cpuregs[10][28] ;
 wire \cpuregs[10][29] ;
 wire \cpuregs[10][2] ;
 wire \cpuregs[10][30] ;
 wire \cpuregs[10][31] ;
 wire \cpuregs[10][3] ;
 wire \cpuregs[10][4] ;
 wire \cpuregs[10][5] ;
 wire \cpuregs[10][6] ;
 wire \cpuregs[10][7] ;
 wire \cpuregs[10][8] ;
 wire \cpuregs[10][9] ;
 wire \cpuregs[11][0] ;
 wire \cpuregs[11][10] ;
 wire \cpuregs[11][11] ;
 wire \cpuregs[11][12] ;
 wire \cpuregs[11][13] ;
 wire \cpuregs[11][14] ;
 wire \cpuregs[11][15] ;
 wire \cpuregs[11][16] ;
 wire \cpuregs[11][17] ;
 wire \cpuregs[11][18] ;
 wire \cpuregs[11][19] ;
 wire \cpuregs[11][1] ;
 wire \cpuregs[11][20] ;
 wire \cpuregs[11][21] ;
 wire \cpuregs[11][22] ;
 wire \cpuregs[11][23] ;
 wire \cpuregs[11][24] ;
 wire \cpuregs[11][25] ;
 wire \cpuregs[11][26] ;
 wire \cpuregs[11][27] ;
 wire \cpuregs[11][28] ;
 wire \cpuregs[11][29] ;
 wire \cpuregs[11][2] ;
 wire \cpuregs[11][30] ;
 wire \cpuregs[11][31] ;
 wire \cpuregs[11][3] ;
 wire \cpuregs[11][4] ;
 wire \cpuregs[11][5] ;
 wire \cpuregs[11][6] ;
 wire \cpuregs[11][7] ;
 wire \cpuregs[11][8] ;
 wire \cpuregs[11][9] ;
 wire \cpuregs[12][0] ;
 wire \cpuregs[12][10] ;
 wire \cpuregs[12][11] ;
 wire \cpuregs[12][12] ;
 wire \cpuregs[12][13] ;
 wire \cpuregs[12][14] ;
 wire \cpuregs[12][15] ;
 wire \cpuregs[12][16] ;
 wire \cpuregs[12][17] ;
 wire \cpuregs[12][18] ;
 wire \cpuregs[12][19] ;
 wire \cpuregs[12][1] ;
 wire \cpuregs[12][20] ;
 wire \cpuregs[12][21] ;
 wire \cpuregs[12][22] ;
 wire \cpuregs[12][23] ;
 wire \cpuregs[12][24] ;
 wire \cpuregs[12][25] ;
 wire \cpuregs[12][26] ;
 wire \cpuregs[12][27] ;
 wire \cpuregs[12][28] ;
 wire \cpuregs[12][29] ;
 wire \cpuregs[12][2] ;
 wire \cpuregs[12][30] ;
 wire \cpuregs[12][31] ;
 wire \cpuregs[12][3] ;
 wire \cpuregs[12][4] ;
 wire \cpuregs[12][5] ;
 wire \cpuregs[12][6] ;
 wire \cpuregs[12][7] ;
 wire \cpuregs[12][8] ;
 wire \cpuregs[12][9] ;
 wire \cpuregs[13][0] ;
 wire \cpuregs[13][10] ;
 wire \cpuregs[13][11] ;
 wire \cpuregs[13][12] ;
 wire \cpuregs[13][13] ;
 wire \cpuregs[13][14] ;
 wire \cpuregs[13][15] ;
 wire \cpuregs[13][16] ;
 wire \cpuregs[13][17] ;
 wire \cpuregs[13][18] ;
 wire \cpuregs[13][19] ;
 wire \cpuregs[13][1] ;
 wire \cpuregs[13][20] ;
 wire \cpuregs[13][21] ;
 wire \cpuregs[13][22] ;
 wire \cpuregs[13][23] ;
 wire \cpuregs[13][24] ;
 wire \cpuregs[13][25] ;
 wire \cpuregs[13][26] ;
 wire \cpuregs[13][27] ;
 wire \cpuregs[13][28] ;
 wire \cpuregs[13][29] ;
 wire \cpuregs[13][2] ;
 wire \cpuregs[13][30] ;
 wire \cpuregs[13][31] ;
 wire \cpuregs[13][3] ;
 wire \cpuregs[13][4] ;
 wire \cpuregs[13][5] ;
 wire \cpuregs[13][6] ;
 wire \cpuregs[13][7] ;
 wire \cpuregs[13][8] ;
 wire \cpuregs[13][9] ;
 wire \cpuregs[14][0] ;
 wire \cpuregs[14][10] ;
 wire \cpuregs[14][11] ;
 wire \cpuregs[14][12] ;
 wire \cpuregs[14][13] ;
 wire \cpuregs[14][14] ;
 wire \cpuregs[14][15] ;
 wire \cpuregs[14][16] ;
 wire \cpuregs[14][17] ;
 wire \cpuregs[14][18] ;
 wire \cpuregs[14][19] ;
 wire \cpuregs[14][1] ;
 wire \cpuregs[14][20] ;
 wire \cpuregs[14][21] ;
 wire \cpuregs[14][22] ;
 wire \cpuregs[14][23] ;
 wire \cpuregs[14][24] ;
 wire \cpuregs[14][25] ;
 wire \cpuregs[14][26] ;
 wire \cpuregs[14][27] ;
 wire \cpuregs[14][28] ;
 wire \cpuregs[14][29] ;
 wire \cpuregs[14][2] ;
 wire \cpuregs[14][30] ;
 wire \cpuregs[14][31] ;
 wire \cpuregs[14][3] ;
 wire \cpuregs[14][4] ;
 wire \cpuregs[14][5] ;
 wire \cpuregs[14][6] ;
 wire \cpuregs[14][7] ;
 wire \cpuregs[14][8] ;
 wire \cpuregs[14][9] ;
 wire \cpuregs[15][0] ;
 wire \cpuregs[15][10] ;
 wire \cpuregs[15][11] ;
 wire \cpuregs[15][12] ;
 wire \cpuregs[15][13] ;
 wire \cpuregs[15][14] ;
 wire \cpuregs[15][15] ;
 wire \cpuregs[15][16] ;
 wire \cpuregs[15][17] ;
 wire \cpuregs[15][18] ;
 wire \cpuregs[15][19] ;
 wire \cpuregs[15][1] ;
 wire \cpuregs[15][20] ;
 wire \cpuregs[15][21] ;
 wire \cpuregs[15][22] ;
 wire \cpuregs[15][23] ;
 wire \cpuregs[15][24] ;
 wire \cpuregs[15][25] ;
 wire \cpuregs[15][26] ;
 wire \cpuregs[15][27] ;
 wire \cpuregs[15][28] ;
 wire \cpuregs[15][29] ;
 wire \cpuregs[15][2] ;
 wire \cpuregs[15][30] ;
 wire \cpuregs[15][31] ;
 wire \cpuregs[15][3] ;
 wire \cpuregs[15][4] ;
 wire \cpuregs[15][5] ;
 wire \cpuregs[15][6] ;
 wire \cpuregs[15][7] ;
 wire \cpuregs[15][8] ;
 wire \cpuregs[15][9] ;
 wire \cpuregs[16][0] ;
 wire \cpuregs[16][10] ;
 wire \cpuregs[16][11] ;
 wire \cpuregs[16][12] ;
 wire \cpuregs[16][13] ;
 wire \cpuregs[16][14] ;
 wire \cpuregs[16][15] ;
 wire \cpuregs[16][16] ;
 wire \cpuregs[16][17] ;
 wire \cpuregs[16][18] ;
 wire \cpuregs[16][19] ;
 wire \cpuregs[16][1] ;
 wire \cpuregs[16][20] ;
 wire \cpuregs[16][21] ;
 wire \cpuregs[16][22] ;
 wire \cpuregs[16][23] ;
 wire \cpuregs[16][24] ;
 wire \cpuregs[16][25] ;
 wire \cpuregs[16][26] ;
 wire \cpuregs[16][27] ;
 wire \cpuregs[16][28] ;
 wire \cpuregs[16][29] ;
 wire \cpuregs[16][2] ;
 wire \cpuregs[16][30] ;
 wire \cpuregs[16][31] ;
 wire \cpuregs[16][3] ;
 wire \cpuregs[16][4] ;
 wire \cpuregs[16][5] ;
 wire \cpuregs[16][6] ;
 wire \cpuregs[16][7] ;
 wire \cpuregs[16][8] ;
 wire \cpuregs[16][9] ;
 wire \cpuregs[17][0] ;
 wire \cpuregs[17][10] ;
 wire \cpuregs[17][11] ;
 wire \cpuregs[17][12] ;
 wire \cpuregs[17][13] ;
 wire \cpuregs[17][14] ;
 wire \cpuregs[17][15] ;
 wire \cpuregs[17][16] ;
 wire \cpuregs[17][17] ;
 wire \cpuregs[17][18] ;
 wire \cpuregs[17][19] ;
 wire \cpuregs[17][1] ;
 wire \cpuregs[17][20] ;
 wire \cpuregs[17][21] ;
 wire \cpuregs[17][22] ;
 wire \cpuregs[17][23] ;
 wire \cpuregs[17][24] ;
 wire \cpuregs[17][25] ;
 wire \cpuregs[17][26] ;
 wire \cpuregs[17][27] ;
 wire \cpuregs[17][28] ;
 wire \cpuregs[17][29] ;
 wire \cpuregs[17][2] ;
 wire \cpuregs[17][30] ;
 wire \cpuregs[17][31] ;
 wire \cpuregs[17][3] ;
 wire \cpuregs[17][4] ;
 wire \cpuregs[17][5] ;
 wire \cpuregs[17][6] ;
 wire \cpuregs[17][7] ;
 wire \cpuregs[17][8] ;
 wire \cpuregs[17][9] ;
 wire \cpuregs[18][0] ;
 wire \cpuregs[18][10] ;
 wire \cpuregs[18][11] ;
 wire \cpuregs[18][12] ;
 wire \cpuregs[18][13] ;
 wire \cpuregs[18][14] ;
 wire \cpuregs[18][15] ;
 wire \cpuregs[18][16] ;
 wire \cpuregs[18][17] ;
 wire \cpuregs[18][18] ;
 wire \cpuregs[18][19] ;
 wire \cpuregs[18][1] ;
 wire \cpuregs[18][20] ;
 wire \cpuregs[18][21] ;
 wire \cpuregs[18][22] ;
 wire \cpuregs[18][23] ;
 wire \cpuregs[18][24] ;
 wire \cpuregs[18][25] ;
 wire \cpuregs[18][26] ;
 wire \cpuregs[18][27] ;
 wire \cpuregs[18][28] ;
 wire \cpuregs[18][29] ;
 wire \cpuregs[18][2] ;
 wire \cpuregs[18][30] ;
 wire \cpuregs[18][31] ;
 wire \cpuregs[18][3] ;
 wire \cpuregs[18][4] ;
 wire \cpuregs[18][5] ;
 wire \cpuregs[18][6] ;
 wire \cpuregs[18][7] ;
 wire \cpuregs[18][8] ;
 wire \cpuregs[18][9] ;
 wire \cpuregs[19][0] ;
 wire \cpuregs[19][10] ;
 wire \cpuregs[19][11] ;
 wire \cpuregs[19][12] ;
 wire \cpuregs[19][13] ;
 wire \cpuregs[19][14] ;
 wire \cpuregs[19][15] ;
 wire \cpuregs[19][16] ;
 wire \cpuregs[19][17] ;
 wire \cpuregs[19][18] ;
 wire \cpuregs[19][19] ;
 wire \cpuregs[19][1] ;
 wire \cpuregs[19][20] ;
 wire \cpuregs[19][21] ;
 wire \cpuregs[19][22] ;
 wire \cpuregs[19][23] ;
 wire \cpuregs[19][24] ;
 wire \cpuregs[19][25] ;
 wire \cpuregs[19][26] ;
 wire \cpuregs[19][27] ;
 wire \cpuregs[19][28] ;
 wire \cpuregs[19][29] ;
 wire \cpuregs[19][2] ;
 wire \cpuregs[19][30] ;
 wire \cpuregs[19][31] ;
 wire \cpuregs[19][3] ;
 wire \cpuregs[19][4] ;
 wire \cpuregs[19][5] ;
 wire \cpuregs[19][6] ;
 wire \cpuregs[19][7] ;
 wire \cpuregs[19][8] ;
 wire \cpuregs[19][9] ;
 wire \cpuregs[1][0] ;
 wire \cpuregs[1][10] ;
 wire \cpuregs[1][11] ;
 wire \cpuregs[1][12] ;
 wire \cpuregs[1][13] ;
 wire \cpuregs[1][14] ;
 wire \cpuregs[1][15] ;
 wire \cpuregs[1][16] ;
 wire \cpuregs[1][17] ;
 wire \cpuregs[1][18] ;
 wire \cpuregs[1][19] ;
 wire \cpuregs[1][1] ;
 wire \cpuregs[1][20] ;
 wire \cpuregs[1][21] ;
 wire \cpuregs[1][22] ;
 wire \cpuregs[1][23] ;
 wire \cpuregs[1][24] ;
 wire \cpuregs[1][25] ;
 wire \cpuregs[1][26] ;
 wire \cpuregs[1][27] ;
 wire \cpuregs[1][28] ;
 wire \cpuregs[1][29] ;
 wire \cpuregs[1][2] ;
 wire \cpuregs[1][30] ;
 wire \cpuregs[1][31] ;
 wire \cpuregs[1][3] ;
 wire \cpuregs[1][4] ;
 wire \cpuregs[1][5] ;
 wire \cpuregs[1][6] ;
 wire \cpuregs[1][7] ;
 wire \cpuregs[1][8] ;
 wire \cpuregs[1][9] ;
 wire \cpuregs[2][0] ;
 wire \cpuregs[2][10] ;
 wire \cpuregs[2][11] ;
 wire \cpuregs[2][12] ;
 wire \cpuregs[2][13] ;
 wire \cpuregs[2][14] ;
 wire \cpuregs[2][15] ;
 wire \cpuregs[2][16] ;
 wire \cpuregs[2][17] ;
 wire \cpuregs[2][18] ;
 wire \cpuregs[2][19] ;
 wire \cpuregs[2][1] ;
 wire \cpuregs[2][20] ;
 wire \cpuregs[2][21] ;
 wire \cpuregs[2][22] ;
 wire \cpuregs[2][23] ;
 wire \cpuregs[2][24] ;
 wire \cpuregs[2][25] ;
 wire \cpuregs[2][26] ;
 wire \cpuregs[2][27] ;
 wire \cpuregs[2][28] ;
 wire \cpuregs[2][29] ;
 wire \cpuregs[2][2] ;
 wire \cpuregs[2][30] ;
 wire \cpuregs[2][31] ;
 wire \cpuregs[2][3] ;
 wire \cpuregs[2][4] ;
 wire \cpuregs[2][5] ;
 wire \cpuregs[2][6] ;
 wire \cpuregs[2][7] ;
 wire \cpuregs[2][8] ;
 wire \cpuregs[2][9] ;
 wire \cpuregs[3][0] ;
 wire \cpuregs[3][10] ;
 wire \cpuregs[3][11] ;
 wire \cpuregs[3][12] ;
 wire \cpuregs[3][13] ;
 wire \cpuregs[3][14] ;
 wire \cpuregs[3][15] ;
 wire \cpuregs[3][16] ;
 wire \cpuregs[3][17] ;
 wire \cpuregs[3][18] ;
 wire \cpuregs[3][19] ;
 wire \cpuregs[3][1] ;
 wire \cpuregs[3][20] ;
 wire \cpuregs[3][21] ;
 wire \cpuregs[3][22] ;
 wire \cpuregs[3][23] ;
 wire \cpuregs[3][24] ;
 wire \cpuregs[3][25] ;
 wire \cpuregs[3][26] ;
 wire \cpuregs[3][27] ;
 wire \cpuregs[3][28] ;
 wire \cpuregs[3][29] ;
 wire \cpuregs[3][2] ;
 wire \cpuregs[3][30] ;
 wire \cpuregs[3][31] ;
 wire \cpuregs[3][3] ;
 wire \cpuregs[3][4] ;
 wire \cpuregs[3][5] ;
 wire \cpuregs[3][6] ;
 wire \cpuregs[3][7] ;
 wire \cpuregs[3][8] ;
 wire \cpuregs[3][9] ;
 wire \cpuregs[4][0] ;
 wire \cpuregs[4][10] ;
 wire \cpuregs[4][11] ;
 wire \cpuregs[4][12] ;
 wire \cpuregs[4][13] ;
 wire \cpuregs[4][14] ;
 wire \cpuregs[4][15] ;
 wire \cpuregs[4][16] ;
 wire \cpuregs[4][17] ;
 wire \cpuregs[4][18] ;
 wire \cpuregs[4][19] ;
 wire \cpuregs[4][1] ;
 wire \cpuregs[4][20] ;
 wire \cpuregs[4][21] ;
 wire \cpuregs[4][22] ;
 wire \cpuregs[4][23] ;
 wire \cpuregs[4][24] ;
 wire \cpuregs[4][25] ;
 wire \cpuregs[4][26] ;
 wire \cpuregs[4][27] ;
 wire \cpuregs[4][28] ;
 wire \cpuregs[4][29] ;
 wire \cpuregs[4][2] ;
 wire \cpuregs[4][30] ;
 wire \cpuregs[4][31] ;
 wire \cpuregs[4][3] ;
 wire \cpuregs[4][4] ;
 wire \cpuregs[4][5] ;
 wire \cpuregs[4][6] ;
 wire \cpuregs[4][7] ;
 wire \cpuregs[4][8] ;
 wire \cpuregs[4][9] ;
 wire \cpuregs[5][0] ;
 wire \cpuregs[5][10] ;
 wire \cpuregs[5][11] ;
 wire \cpuregs[5][12] ;
 wire \cpuregs[5][13] ;
 wire \cpuregs[5][14] ;
 wire \cpuregs[5][15] ;
 wire \cpuregs[5][16] ;
 wire \cpuregs[5][17] ;
 wire \cpuregs[5][18] ;
 wire \cpuregs[5][19] ;
 wire \cpuregs[5][1] ;
 wire \cpuregs[5][20] ;
 wire \cpuregs[5][21] ;
 wire \cpuregs[5][22] ;
 wire \cpuregs[5][23] ;
 wire \cpuregs[5][24] ;
 wire \cpuregs[5][25] ;
 wire \cpuregs[5][26] ;
 wire \cpuregs[5][27] ;
 wire \cpuregs[5][28] ;
 wire \cpuregs[5][29] ;
 wire \cpuregs[5][2] ;
 wire \cpuregs[5][30] ;
 wire \cpuregs[5][31] ;
 wire \cpuregs[5][3] ;
 wire \cpuregs[5][4] ;
 wire \cpuregs[5][5] ;
 wire \cpuregs[5][6] ;
 wire \cpuregs[5][7] ;
 wire \cpuregs[5][8] ;
 wire \cpuregs[5][9] ;
 wire \cpuregs[6][0] ;
 wire \cpuregs[6][10] ;
 wire \cpuregs[6][11] ;
 wire \cpuregs[6][12] ;
 wire \cpuregs[6][13] ;
 wire \cpuregs[6][14] ;
 wire \cpuregs[6][15] ;
 wire \cpuregs[6][16] ;
 wire \cpuregs[6][17] ;
 wire \cpuregs[6][18] ;
 wire \cpuregs[6][19] ;
 wire \cpuregs[6][1] ;
 wire \cpuregs[6][20] ;
 wire \cpuregs[6][21] ;
 wire \cpuregs[6][22] ;
 wire \cpuregs[6][23] ;
 wire \cpuregs[6][24] ;
 wire \cpuregs[6][25] ;
 wire \cpuregs[6][26] ;
 wire \cpuregs[6][27] ;
 wire \cpuregs[6][28] ;
 wire \cpuregs[6][29] ;
 wire \cpuregs[6][2] ;
 wire \cpuregs[6][30] ;
 wire \cpuregs[6][31] ;
 wire \cpuregs[6][3] ;
 wire \cpuregs[6][4] ;
 wire \cpuregs[6][5] ;
 wire \cpuregs[6][6] ;
 wire \cpuregs[6][7] ;
 wire \cpuregs[6][8] ;
 wire \cpuregs[6][9] ;
 wire \cpuregs[7][0] ;
 wire \cpuregs[7][10] ;
 wire \cpuregs[7][11] ;
 wire \cpuregs[7][12] ;
 wire \cpuregs[7][13] ;
 wire \cpuregs[7][14] ;
 wire \cpuregs[7][15] ;
 wire \cpuregs[7][16] ;
 wire \cpuregs[7][17] ;
 wire \cpuregs[7][18] ;
 wire \cpuregs[7][19] ;
 wire \cpuregs[7][1] ;
 wire \cpuregs[7][20] ;
 wire \cpuregs[7][21] ;
 wire \cpuregs[7][22] ;
 wire \cpuregs[7][23] ;
 wire \cpuregs[7][24] ;
 wire \cpuregs[7][25] ;
 wire \cpuregs[7][26] ;
 wire \cpuregs[7][27] ;
 wire \cpuregs[7][28] ;
 wire \cpuregs[7][29] ;
 wire \cpuregs[7][2] ;
 wire \cpuregs[7][30] ;
 wire \cpuregs[7][31] ;
 wire \cpuregs[7][3] ;
 wire \cpuregs[7][4] ;
 wire \cpuregs[7][5] ;
 wire \cpuregs[7][6] ;
 wire \cpuregs[7][7] ;
 wire \cpuregs[7][8] ;
 wire \cpuregs[7][9] ;
 wire \cpuregs[8][0] ;
 wire \cpuregs[8][10] ;
 wire \cpuregs[8][11] ;
 wire \cpuregs[8][12] ;
 wire \cpuregs[8][13] ;
 wire \cpuregs[8][14] ;
 wire \cpuregs[8][15] ;
 wire \cpuregs[8][16] ;
 wire \cpuregs[8][17] ;
 wire \cpuregs[8][18] ;
 wire \cpuregs[8][19] ;
 wire \cpuregs[8][1] ;
 wire \cpuregs[8][20] ;
 wire \cpuregs[8][21] ;
 wire \cpuregs[8][22] ;
 wire \cpuregs[8][23] ;
 wire \cpuregs[8][24] ;
 wire \cpuregs[8][25] ;
 wire \cpuregs[8][26] ;
 wire \cpuregs[8][27] ;
 wire \cpuregs[8][28] ;
 wire \cpuregs[8][29] ;
 wire \cpuregs[8][2] ;
 wire \cpuregs[8][30] ;
 wire \cpuregs[8][31] ;
 wire \cpuregs[8][3] ;
 wire \cpuregs[8][4] ;
 wire \cpuregs[8][5] ;
 wire \cpuregs[8][6] ;
 wire \cpuregs[8][7] ;
 wire \cpuregs[8][8] ;
 wire \cpuregs[8][9] ;
 wire \cpuregs[9][0] ;
 wire \cpuregs[9][10] ;
 wire \cpuregs[9][11] ;
 wire \cpuregs[9][12] ;
 wire \cpuregs[9][13] ;
 wire \cpuregs[9][14] ;
 wire \cpuregs[9][15] ;
 wire \cpuregs[9][16] ;
 wire \cpuregs[9][17] ;
 wire \cpuregs[9][18] ;
 wire \cpuregs[9][19] ;
 wire \cpuregs[9][1] ;
 wire \cpuregs[9][20] ;
 wire \cpuregs[9][21] ;
 wire \cpuregs[9][22] ;
 wire \cpuregs[9][23] ;
 wire \cpuregs[9][24] ;
 wire \cpuregs[9][25] ;
 wire \cpuregs[9][26] ;
 wire \cpuregs[9][27] ;
 wire \cpuregs[9][28] ;
 wire \cpuregs[9][29] ;
 wire \cpuregs[9][2] ;
 wire \cpuregs[9][30] ;
 wire \cpuregs[9][31] ;
 wire \cpuregs[9][3] ;
 wire \cpuregs[9][4] ;
 wire \cpuregs[9][5] ;
 wire \cpuregs[9][6] ;
 wire \cpuregs[9][7] ;
 wire \cpuregs[9][8] ;
 wire \cpuregs[9][9] ;
 wire \cpuregs_rs1[0] ;
 wire \cpuregs_rs1[10] ;
 wire \cpuregs_rs1[11] ;
 wire \cpuregs_rs1[12] ;
 wire \cpuregs_rs1[13] ;
 wire \cpuregs_rs1[14] ;
 wire \cpuregs_rs1[15] ;
 wire \cpuregs_rs1[16] ;
 wire \cpuregs_rs1[17] ;
 wire \cpuregs_rs1[18] ;
 wire \cpuregs_rs1[19] ;
 wire \cpuregs_rs1[1] ;
 wire \cpuregs_rs1[20] ;
 wire \cpuregs_rs1[21] ;
 wire \cpuregs_rs1[22] ;
 wire \cpuregs_rs1[23] ;
 wire \cpuregs_rs1[24] ;
 wire \cpuregs_rs1[25] ;
 wire \cpuregs_rs1[26] ;
 wire \cpuregs_rs1[27] ;
 wire \cpuregs_rs1[28] ;
 wire \cpuregs_rs1[29] ;
 wire \cpuregs_rs1[2] ;
 wire \cpuregs_rs1[30] ;
 wire \cpuregs_rs1[31] ;
 wire \cpuregs_rs1[3] ;
 wire \cpuregs_rs1[4] ;
 wire \cpuregs_rs1[5] ;
 wire \cpuregs_rs1[6] ;
 wire \cpuregs_rs1[7] ;
 wire \cpuregs_rs1[8] ;
 wire \cpuregs_rs1[9] ;
 wire \cpuregs_wrdata[0] ;
 wire \cpuregs_wrdata[10] ;
 wire \cpuregs_wrdata[11] ;
 wire \cpuregs_wrdata[12] ;
 wire \cpuregs_wrdata[13] ;
 wire \cpuregs_wrdata[14] ;
 wire \cpuregs_wrdata[15] ;
 wire \cpuregs_wrdata[16] ;
 wire \cpuregs_wrdata[17] ;
 wire \cpuregs_wrdata[18] ;
 wire \cpuregs_wrdata[19] ;
 wire \cpuregs_wrdata[1] ;
 wire \cpuregs_wrdata[20] ;
 wire \cpuregs_wrdata[21] ;
 wire \cpuregs_wrdata[22] ;
 wire \cpuregs_wrdata[23] ;
 wire \cpuregs_wrdata[24] ;
 wire \cpuregs_wrdata[25] ;
 wire \cpuregs_wrdata[26] ;
 wire \cpuregs_wrdata[27] ;
 wire \cpuregs_wrdata[28] ;
 wire \cpuregs_wrdata[29] ;
 wire \cpuregs_wrdata[2] ;
 wire \cpuregs_wrdata[30] ;
 wire \cpuregs_wrdata[31] ;
 wire \cpuregs_wrdata[3] ;
 wire \cpuregs_wrdata[4] ;
 wire \cpuregs_wrdata[5] ;
 wire \cpuregs_wrdata[6] ;
 wire \cpuregs_wrdata[7] ;
 wire \cpuregs_wrdata[8] ;
 wire \cpuregs_wrdata[9] ;
 wire \decoded_imm[0] ;
 wire \decoded_imm[10] ;
 wire \decoded_imm[11] ;
 wire \decoded_imm[12] ;
 wire \decoded_imm[13] ;
 wire \decoded_imm[14] ;
 wire \decoded_imm[15] ;
 wire \decoded_imm[16] ;
 wire \decoded_imm[17] ;
 wire \decoded_imm[18] ;
 wire \decoded_imm[19] ;
 wire \decoded_imm[1] ;
 wire \decoded_imm[20] ;
 wire \decoded_imm[21] ;
 wire \decoded_imm[22] ;
 wire \decoded_imm[23] ;
 wire \decoded_imm[24] ;
 wire \decoded_imm[25] ;
 wire \decoded_imm[26] ;
 wire \decoded_imm[27] ;
 wire \decoded_imm[28] ;
 wire \decoded_imm[29] ;
 wire \decoded_imm[2] ;
 wire \decoded_imm[30] ;
 wire \decoded_imm[31] ;
 wire \decoded_imm[3] ;
 wire \decoded_imm[4] ;
 wire \decoded_imm[5] ;
 wire \decoded_imm[6] ;
 wire \decoded_imm[7] ;
 wire \decoded_imm[8] ;
 wire \decoded_imm[9] ;
 wire \decoded_imm_uj[10] ;
 wire \decoded_imm_uj[11] ;
 wire \decoded_imm_uj[12] ;
 wire \decoded_imm_uj[13] ;
 wire \decoded_imm_uj[14] ;
 wire \decoded_imm_uj[15] ;
 wire \decoded_imm_uj[16] ;
 wire \decoded_imm_uj[17] ;
 wire \decoded_imm_uj[18] ;
 wire \decoded_imm_uj[19] ;
 wire \decoded_imm_uj[1] ;
 wire \decoded_imm_uj[20] ;
 wire \decoded_imm_uj[2] ;
 wire \decoded_imm_uj[3] ;
 wire \decoded_imm_uj[4] ;
 wire \decoded_imm_uj[5] ;
 wire \decoded_imm_uj[6] ;
 wire \decoded_imm_uj[7] ;
 wire \decoded_imm_uj[8] ;
 wire \decoded_imm_uj[9] ;
 wire \decoded_rd[0] ;
 wire \decoded_rd[1] ;
 wire \decoded_rd[2] ;
 wire \decoded_rd[3] ;
 wire \decoded_rd[4] ;
 wire \decoded_rs1[0] ;
 wire \decoded_rs1[1] ;
 wire \decoded_rs1[2] ;
 wire \decoded_rs1[3] ;
 wire \decoded_rs1[4] ;
 wire decoder_pseudo_trigger;
 wire decoder_trigger;
 wire do_waitirq;
 wire instr_add;
 wire instr_addi;
 wire instr_and;
 wire instr_andi;
 wire instr_auipc;
 wire instr_beq;
 wire instr_bge;
 wire instr_bgeu;
 wire instr_blt;
 wire instr_bltu;
 wire instr_bne;
 wire instr_ecall_ebreak;
 wire instr_getq;
 wire instr_jal;
 wire instr_jalr;
 wire instr_lb;
 wire instr_lbu;
 wire instr_lh;
 wire instr_lhu;
 wire instr_lui;
 wire instr_lw;
 wire instr_maskirq;
 wire instr_or;
 wire instr_ori;
 wire instr_rdcycle;
 wire instr_rdcycleh;
 wire instr_rdinstr;
 wire instr_rdinstrh;
 wire instr_retirq;
 wire instr_sb;
 wire instr_setq;
 wire instr_sh;
 wire instr_sll;
 wire instr_slli;
 wire instr_slt;
 wire instr_slti;
 wire instr_sltiu;
 wire instr_sltu;
 wire instr_sra;
 wire instr_srai;
 wire instr_srl;
 wire instr_srli;
 wire instr_sub;
 wire instr_sw;
 wire instr_timer;
 wire instr_waitirq;
 wire instr_xor;
 wire instr_xori;
 wire irq_active;
 wire irq_delay;
 wire \irq_mask[0] ;
 wire \irq_mask[10] ;
 wire \irq_mask[11] ;
 wire \irq_mask[12] ;
 wire \irq_mask[13] ;
 wire \irq_mask[14] ;
 wire \irq_mask[15] ;
 wire \irq_mask[16] ;
 wire \irq_mask[17] ;
 wire \irq_mask[18] ;
 wire \irq_mask[19] ;
 wire \irq_mask[1] ;
 wire \irq_mask[20] ;
 wire \irq_mask[21] ;
 wire \irq_mask[22] ;
 wire \irq_mask[23] ;
 wire \irq_mask[24] ;
 wire \irq_mask[25] ;
 wire \irq_mask[26] ;
 wire \irq_mask[27] ;
 wire \irq_mask[28] ;
 wire \irq_mask[29] ;
 wire \irq_mask[2] ;
 wire \irq_mask[30] ;
 wire \irq_mask[31] ;
 wire \irq_mask[3] ;
 wire \irq_mask[4] ;
 wire \irq_mask[5] ;
 wire \irq_mask[6] ;
 wire \irq_mask[7] ;
 wire \irq_mask[8] ;
 wire \irq_mask[9] ;
 wire \irq_pending[0] ;
 wire \irq_pending[10] ;
 wire \irq_pending[11] ;
 wire \irq_pending[12] ;
 wire \irq_pending[13] ;
 wire \irq_pending[14] ;
 wire \irq_pending[15] ;
 wire \irq_pending[16] ;
 wire \irq_pending[17] ;
 wire \irq_pending[18] ;
 wire \irq_pending[19] ;
 wire \irq_pending[1] ;
 wire \irq_pending[20] ;
 wire \irq_pending[21] ;
 wire \irq_pending[22] ;
 wire \irq_pending[23] ;
 wire \irq_pending[24] ;
 wire \irq_pending[25] ;
 wire \irq_pending[26] ;
 wire \irq_pending[27] ;
 wire \irq_pending[28] ;
 wire \irq_pending[29] ;
 wire \irq_pending[2] ;
 wire \irq_pending[30] ;
 wire \irq_pending[31] ;
 wire \irq_pending[3] ;
 wire \irq_pending[4] ;
 wire \irq_pending[5] ;
 wire \irq_pending[6] ;
 wire \irq_pending[7] ;
 wire \irq_pending[8] ;
 wire \irq_pending[9] ;
 wire \irq_state[0] ;
 wire \irq_state[1] ;
 wire is_alu_reg_imm;
 wire is_alu_reg_reg;
 wire is_beq_bne_blt_bge_bltu_bgeu;
 wire is_compare;
 wire is_jalr_addi_slti_sltiu_xori_ori_andi;
 wire is_lb_lh_lw_lbu_lhu;
 wire is_lui_auipc_jal;
 wire is_sb_sh_sw;
 wire is_slli_srli_srai;
 wire is_slti_blt_slt;
 wire is_sltiu_bltu_sltu;
 wire latched_branch;
 wire latched_is_lb;
 wire latched_is_lh;
 wire \latched_rd[0] ;
 wire \latched_rd[1] ;
 wire \latched_rd[2] ;
 wire \latched_rd[3] ;
 wire \latched_rd[4] ;
 wire latched_stalu;
 wire latched_store;
 wire mem_do_prefetch;
 wire mem_do_rdata;
 wire mem_do_rinst;
 wire mem_do_wdata;
 wire \mem_rdata_latched[10] ;
 wire \mem_rdata_latched[11] ;
 wire \mem_rdata_latched[12] ;
 wire \mem_rdata_latched[13] ;
 wire \mem_rdata_latched[14] ;
 wire \mem_rdata_latched[15] ;
 wire \mem_rdata_latched[16] ;
 wire \mem_rdata_latched[17] ;
 wire \mem_rdata_latched[18] ;
 wire \mem_rdata_latched[19] ;
 wire \mem_rdata_latched[20] ;
 wire \mem_rdata_latched[21] ;
 wire \mem_rdata_latched[22] ;
 wire \mem_rdata_latched[23] ;
 wire \mem_rdata_latched[24] ;
 wire \mem_rdata_latched[25] ;
 wire \mem_rdata_latched[26] ;
 wire \mem_rdata_latched[27] ;
 wire \mem_rdata_latched[28] ;
 wire \mem_rdata_latched[29] ;
 wire \mem_rdata_latched[30] ;
 wire \mem_rdata_latched[31] ;
 wire \mem_rdata_latched[7] ;
 wire \mem_rdata_latched[8] ;
 wire \mem_rdata_latched[9] ;
 wire \mem_rdata_q[0] ;
 wire \mem_rdata_q[10] ;
 wire \mem_rdata_q[11] ;
 wire \mem_rdata_q[12] ;
 wire \mem_rdata_q[13] ;
 wire \mem_rdata_q[14] ;
 wire \mem_rdata_q[15] ;
 wire \mem_rdata_q[16] ;
 wire \mem_rdata_q[17] ;
 wire \mem_rdata_q[18] ;
 wire \mem_rdata_q[19] ;
 wire \mem_rdata_q[1] ;
 wire \mem_rdata_q[20] ;
 wire \mem_rdata_q[21] ;
 wire \mem_rdata_q[22] ;
 wire \mem_rdata_q[23] ;
 wire \mem_rdata_q[24] ;
 wire \mem_rdata_q[25] ;
 wire \mem_rdata_q[26] ;
 wire \mem_rdata_q[27] ;
 wire \mem_rdata_q[28] ;
 wire \mem_rdata_q[29] ;
 wire \mem_rdata_q[2] ;
 wire \mem_rdata_q[30] ;
 wire \mem_rdata_q[31] ;
 wire \mem_rdata_q[3] ;
 wire \mem_rdata_q[4] ;
 wire \mem_rdata_q[5] ;
 wire \mem_rdata_q[6] ;
 wire \mem_rdata_q[7] ;
 wire \mem_rdata_q[8] ;
 wire \mem_rdata_q[9] ;
 wire \mem_state[0] ;
 wire \mem_state[1] ;
 wire \mem_wordsize[0] ;
 wire \mem_wordsize[1] ;
 wire \mem_wordsize[2] ;
 wire mem_xfer;
 wire \pcpi_mul.active[0] ;
 wire \pcpi_mul.active[1] ;
 wire \pcpi_mul.instr_any_mulh ;
 wire \pcpi_mul.rd[0] ;
 wire \pcpi_mul.rd[10] ;
 wire \pcpi_mul.rd[11] ;
 wire \pcpi_mul.rd[12] ;
 wire \pcpi_mul.rd[13] ;
 wire \pcpi_mul.rd[14] ;
 wire \pcpi_mul.rd[15] ;
 wire \pcpi_mul.rd[16] ;
 wire \pcpi_mul.rd[17] ;
 wire \pcpi_mul.rd[18] ;
 wire \pcpi_mul.rd[19] ;
 wire \pcpi_mul.rd[1] ;
 wire \pcpi_mul.rd[20] ;
 wire \pcpi_mul.rd[21] ;
 wire \pcpi_mul.rd[22] ;
 wire \pcpi_mul.rd[23] ;
 wire \pcpi_mul.rd[24] ;
 wire \pcpi_mul.rd[25] ;
 wire \pcpi_mul.rd[26] ;
 wire \pcpi_mul.rd[27] ;
 wire \pcpi_mul.rd[28] ;
 wire \pcpi_mul.rd[29] ;
 wire \pcpi_mul.rd[2] ;
 wire \pcpi_mul.rd[30] ;
 wire \pcpi_mul.rd[31] ;
 wire \pcpi_mul.rd[32] ;
 wire \pcpi_mul.rd[33] ;
 wire \pcpi_mul.rd[34] ;
 wire \pcpi_mul.rd[35] ;
 wire \pcpi_mul.rd[36] ;
 wire \pcpi_mul.rd[37] ;
 wire \pcpi_mul.rd[38] ;
 wire \pcpi_mul.rd[39] ;
 wire \pcpi_mul.rd[3] ;
 wire \pcpi_mul.rd[40] ;
 wire \pcpi_mul.rd[41] ;
 wire \pcpi_mul.rd[42] ;
 wire \pcpi_mul.rd[43] ;
 wire \pcpi_mul.rd[44] ;
 wire \pcpi_mul.rd[45] ;
 wire \pcpi_mul.rd[46] ;
 wire \pcpi_mul.rd[47] ;
 wire \pcpi_mul.rd[48] ;
 wire \pcpi_mul.rd[49] ;
 wire \pcpi_mul.rd[4] ;
 wire \pcpi_mul.rd[50] ;
 wire \pcpi_mul.rd[51] ;
 wire \pcpi_mul.rd[52] ;
 wire \pcpi_mul.rd[53] ;
 wire \pcpi_mul.rd[54] ;
 wire \pcpi_mul.rd[55] ;
 wire \pcpi_mul.rd[56] ;
 wire \pcpi_mul.rd[57] ;
 wire \pcpi_mul.rd[58] ;
 wire \pcpi_mul.rd[59] ;
 wire \pcpi_mul.rd[5] ;
 wire \pcpi_mul.rd[60] ;
 wire \pcpi_mul.rd[61] ;
 wire \pcpi_mul.rd[62] ;
 wire \pcpi_mul.rd[63] ;
 wire \pcpi_mul.rd[6] ;
 wire \pcpi_mul.rd[7] ;
 wire \pcpi_mul.rd[8] ;
 wire \pcpi_mul.rd[9] ;
 wire \pcpi_mul.rs1[0] ;
 wire \pcpi_mul.rs1[10] ;
 wire \pcpi_mul.rs1[11] ;
 wire \pcpi_mul.rs1[12] ;
 wire \pcpi_mul.rs1[13] ;
 wire \pcpi_mul.rs1[14] ;
 wire \pcpi_mul.rs1[15] ;
 wire \pcpi_mul.rs1[16] ;
 wire \pcpi_mul.rs1[17] ;
 wire \pcpi_mul.rs1[18] ;
 wire \pcpi_mul.rs1[19] ;
 wire \pcpi_mul.rs1[1] ;
 wire \pcpi_mul.rs1[20] ;
 wire \pcpi_mul.rs1[21] ;
 wire \pcpi_mul.rs1[22] ;
 wire \pcpi_mul.rs1[23] ;
 wire \pcpi_mul.rs1[24] ;
 wire \pcpi_mul.rs1[25] ;
 wire \pcpi_mul.rs1[26] ;
 wire \pcpi_mul.rs1[27] ;
 wire \pcpi_mul.rs1[28] ;
 wire \pcpi_mul.rs1[29] ;
 wire \pcpi_mul.rs1[2] ;
 wire \pcpi_mul.rs1[30] ;
 wire \pcpi_mul.rs1[31] ;
 wire \pcpi_mul.rs1[32] ;
 wire \pcpi_mul.rs1[3] ;
 wire \pcpi_mul.rs1[4] ;
 wire \pcpi_mul.rs1[5] ;
 wire \pcpi_mul.rs1[6] ;
 wire \pcpi_mul.rs1[7] ;
 wire \pcpi_mul.rs1[8] ;
 wire \pcpi_mul.rs1[9] ;
 wire \pcpi_mul.rs2[0] ;
 wire \pcpi_mul.rs2[10] ;
 wire \pcpi_mul.rs2[11] ;
 wire \pcpi_mul.rs2[12] ;
 wire \pcpi_mul.rs2[13] ;
 wire \pcpi_mul.rs2[14] ;
 wire \pcpi_mul.rs2[15] ;
 wire \pcpi_mul.rs2[16] ;
 wire \pcpi_mul.rs2[17] ;
 wire \pcpi_mul.rs2[18] ;
 wire \pcpi_mul.rs2[19] ;
 wire \pcpi_mul.rs2[1] ;
 wire \pcpi_mul.rs2[20] ;
 wire \pcpi_mul.rs2[21] ;
 wire \pcpi_mul.rs2[22] ;
 wire \pcpi_mul.rs2[23] ;
 wire \pcpi_mul.rs2[24] ;
 wire \pcpi_mul.rs2[25] ;
 wire \pcpi_mul.rs2[26] ;
 wire \pcpi_mul.rs2[27] ;
 wire \pcpi_mul.rs2[28] ;
 wire \pcpi_mul.rs2[29] ;
 wire \pcpi_mul.rs2[2] ;
 wire \pcpi_mul.rs2[30] ;
 wire \pcpi_mul.rs2[31] ;
 wire \pcpi_mul.rs2[32] ;
 wire \pcpi_mul.rs2[3] ;
 wire \pcpi_mul.rs2[4] ;
 wire \pcpi_mul.rs2[5] ;
 wire \pcpi_mul.rs2[6] ;
 wire \pcpi_mul.rs2[7] ;
 wire \pcpi_mul.rs2[8] ;
 wire \pcpi_mul.rs2[9] ;
 wire \pcpi_mul.shift_out ;
 wire pcpi_timeout;
 wire \pcpi_timeout_counter[0] ;
 wire \pcpi_timeout_counter[1] ;
 wire \pcpi_timeout_counter[2] ;
 wire \pcpi_timeout_counter[3] ;
 wire \reg_next_pc[0] ;
 wire \reg_next_pc[10] ;
 wire \reg_next_pc[11] ;
 wire \reg_next_pc[12] ;
 wire \reg_next_pc[13] ;
 wire \reg_next_pc[14] ;
 wire \reg_next_pc[15] ;
 wire \reg_next_pc[16] ;
 wire \reg_next_pc[17] ;
 wire \reg_next_pc[18] ;
 wire \reg_next_pc[19] ;
 wire \reg_next_pc[1] ;
 wire \reg_next_pc[20] ;
 wire \reg_next_pc[21] ;
 wire \reg_next_pc[22] ;
 wire \reg_next_pc[23] ;
 wire \reg_next_pc[24] ;
 wire \reg_next_pc[25] ;
 wire \reg_next_pc[26] ;
 wire \reg_next_pc[27] ;
 wire \reg_next_pc[28] ;
 wire \reg_next_pc[29] ;
 wire \reg_next_pc[2] ;
 wire \reg_next_pc[30] ;
 wire \reg_next_pc[31] ;
 wire \reg_next_pc[3] ;
 wire \reg_next_pc[4] ;
 wire \reg_next_pc[5] ;
 wire \reg_next_pc[6] ;
 wire \reg_next_pc[7] ;
 wire \reg_next_pc[8] ;
 wire \reg_next_pc[9] ;
 wire \reg_out[0] ;
 wire \reg_out[10] ;
 wire \reg_out[11] ;
 wire \reg_out[12] ;
 wire \reg_out[13] ;
 wire \reg_out[14] ;
 wire \reg_out[15] ;
 wire \reg_out[16] ;
 wire \reg_out[17] ;
 wire \reg_out[18] ;
 wire \reg_out[19] ;
 wire \reg_out[1] ;
 wire \reg_out[20] ;
 wire \reg_out[21] ;
 wire \reg_out[22] ;
 wire \reg_out[23] ;
 wire \reg_out[24] ;
 wire \reg_out[25] ;
 wire \reg_out[26] ;
 wire \reg_out[27] ;
 wire \reg_out[28] ;
 wire \reg_out[29] ;
 wire \reg_out[2] ;
 wire \reg_out[30] ;
 wire \reg_out[31] ;
 wire \reg_out[3] ;
 wire \reg_out[4] ;
 wire \reg_out[5] ;
 wire \reg_out[6] ;
 wire \reg_out[7] ;
 wire \reg_out[8] ;
 wire \reg_out[9] ;
 wire \reg_pc[10] ;
 wire \reg_pc[11] ;
 wire \reg_pc[12] ;
 wire \reg_pc[13] ;
 wire \reg_pc[14] ;
 wire \reg_pc[15] ;
 wire \reg_pc[16] ;
 wire \reg_pc[17] ;
 wire \reg_pc[18] ;
 wire \reg_pc[19] ;
 wire \reg_pc[1] ;
 wire \reg_pc[20] ;
 wire \reg_pc[21] ;
 wire \reg_pc[22] ;
 wire \reg_pc[23] ;
 wire \reg_pc[24] ;
 wire \reg_pc[25] ;
 wire \reg_pc[26] ;
 wire \reg_pc[27] ;
 wire \reg_pc[28] ;
 wire \reg_pc[29] ;
 wire \reg_pc[2] ;
 wire \reg_pc[30] ;
 wire \reg_pc[31] ;
 wire \reg_pc[3] ;
 wire \reg_pc[4] ;
 wire \reg_pc[5] ;
 wire \reg_pc[6] ;
 wire \reg_pc[7] ;
 wire \reg_pc[8] ;
 wire \reg_pc[9] ;
 wire \timer[0] ;
 wire \timer[10] ;
 wire \timer[11] ;
 wire \timer[12] ;
 wire \timer[13] ;
 wire \timer[14] ;
 wire \timer[15] ;
 wire \timer[16] ;
 wire \timer[17] ;
 wire \timer[18] ;
 wire \timer[19] ;
 wire \timer[1] ;
 wire \timer[20] ;
 wire \timer[21] ;
 wire \timer[22] ;
 wire \timer[23] ;
 wire \timer[24] ;
 wire \timer[25] ;
 wire \timer[26] ;
 wire \timer[27] ;
 wire \timer[28] ;
 wire \timer[29] ;
 wire \timer[2] ;
 wire \timer[30] ;
 wire \timer[31] ;
 wire \timer[3] ;
 wire \timer[4] ;
 wire \timer[5] ;
 wire \timer[6] ;
 wire \timer[7] ;
 wire \timer[8] ;
 wire \timer[9] ;

 sky130_fd_sc_hd__buf_1 _13031_ (.A(resetn),
    .X(_10443_));
 sky130_fd_sc_hd__buf_1 _13032_ (.A(_10443_),
    .X(_10444_));
 sky130_fd_sc_hd__nand2_2 _13033_ (.A(mem_valid),
    .B(mem_ready),
    .Y(_10445_));
 sky130_vsdinv _13034_ (.A(_10445_),
    .Y(_10446_));
 sky130_fd_sc_hd__buf_1 _13035_ (.A(_10446_),
    .X(_10447_));
 sky130_vsdinv _13036_ (.A(\mem_state[1] ),
    .Y(_10448_));
 sky130_vsdinv _13037_ (.A(\mem_state[0] ),
    .Y(_10449_));
 sky130_fd_sc_hd__nor2_2 _13038_ (.A(_10448_),
    .B(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__o21a_2 _13039_ (.A1(mem_do_wdata),
    .A2(mem_do_rdata),
    .B1(_10446_),
    .X(_10451_));
 sky130_fd_sc_hd__or2_2 _13040_ (.A(\mem_state[1] ),
    .B(\mem_state[0] ),
    .X(_10452_));
 sky130_fd_sc_hd__o221a_2 _13041_ (.A1(_10447_),
    .A2(_10450_),
    .B1(mem_do_rinst),
    .B2(_10451_),
    .C1(_10452_),
    .X(_10453_));
 sky130_fd_sc_hd__nand2_2 _13042_ (.A(resetn),
    .B(_10453_),
    .Y(_10454_));
 sky130_fd_sc_hd__nand2_2 _13043_ (.A(mem_do_prefetch),
    .B(_10454_),
    .Y(_10455_));
 sky130_vsdinv _13044_ (.A(mem_do_rdata),
    .Y(_10456_));
 sky130_fd_sc_hd__buf_1 _13045_ (.A(\cpu_state[6] ),
    .X(_10457_));
 sky130_vsdinv _13046_ (.A(_10457_),
    .Y(_10458_));
 sky130_fd_sc_hd__buf_1 _13047_ (.A(_10458_),
    .X(_10459_));
 sky130_fd_sc_hd__nor2_2 _13048_ (.A(_10456_),
    .B(_10459_),
    .Y(_00319_));
 sky130_fd_sc_hd__a31o_2 _13049_ (.A1(_10444_),
    .A2(_10455_),
    .A3(_00319_),
    .B1(_00332_),
    .X(_10460_));
 sky130_vsdinv _13050_ (.A(_10460_),
    .Y(_10461_));
 sky130_fd_sc_hd__and2_2 _13051_ (.A(instr_lb),
    .B(_10457_),
    .X(_10462_));
 sky130_fd_sc_hd__buf_1 _13052_ (.A(_10443_),
    .X(_10463_));
 sky130_fd_sc_hd__buf_1 _13053_ (.A(_10463_),
    .X(_10464_));
 sky130_fd_sc_hd__o221a_2 _13054_ (.A1(latched_is_lb),
    .A2(_10461_),
    .B1(_10460_),
    .B2(_10462_),
    .C1(_10464_),
    .X(_04071_));
 sky130_fd_sc_hd__and2_2 _13055_ (.A(instr_lh),
    .B(_10457_),
    .X(_10465_));
 sky130_fd_sc_hd__buf_1 _13056_ (.A(_10444_),
    .X(_10466_));
 sky130_fd_sc_hd__buf_1 _13057_ (.A(_10466_),
    .X(_10467_));
 sky130_fd_sc_hd__o221a_2 _13058_ (.A1(latched_is_lh),
    .A2(_10461_),
    .B1(_10460_),
    .B2(_10465_),
    .C1(_10467_),
    .X(_04070_));
 sky130_vsdinv _13059_ (.A(\cpu_state[2] ),
    .Y(_10468_));
 sky130_fd_sc_hd__buf_1 _13060_ (.A(_10468_),
    .X(_10469_));
 sky130_fd_sc_hd__buf_1 _13061_ (.A(_10469_),
    .X(_10470_));
 sky130_fd_sc_hd__o21ba_2 _13062_ (.A1(instr_retirq),
    .A2(_10470_),
    .B1_N(_00331_),
    .X(_10471_));
 sky130_vsdinv _13063_ (.A(_10471_),
    .Y(_10472_));
 sky130_fd_sc_hd__buf_1 _13064_ (.A(latched_branch),
    .X(_10473_));
 sky130_fd_sc_hd__o221a_2 _13065_ (.A1(_12980_),
    .A2(_10472_),
    .B1(_10473_),
    .B2(_10471_),
    .C1(_10467_),
    .X(_04069_));
 sky130_vsdinv _13066_ (.A(resetn),
    .Y(_10474_));
 sky130_fd_sc_hd__buf_1 _13067_ (.A(_10474_),
    .X(_10475_));
 sky130_fd_sc_hd__buf_1 _13068_ (.A(_10475_),
    .X(_10476_));
 sky130_fd_sc_hd__buf_1 _13069_ (.A(_10476_),
    .X(_10477_));
 sky130_fd_sc_hd__or2_2 _13070_ (.A(_10477_),
    .B(trap),
    .X(_10478_));
 sky130_vsdinv _13071_ (.A(_10478_),
    .Y(_10479_));
 sky130_fd_sc_hd__buf_1 _13072_ (.A(_10479_),
    .X(_10480_));
 sky130_fd_sc_hd__buf_1 _13073_ (.A(_10477_),
    .X(_10481_));
 sky130_fd_sc_hd__buf_1 _13074_ (.A(_10481_),
    .X(_10482_));
 sky130_fd_sc_hd__or2_2 _13075_ (.A(mem_do_rinst),
    .B(mem_do_prefetch),
    .X(_10483_));
 sky130_fd_sc_hd__or2_2 _13076_ (.A(mem_do_rdata),
    .B(_10483_),
    .X(_10484_));
 sky130_vsdinv _13077_ (.A(trap),
    .Y(_10485_));
 sky130_fd_sc_hd__a221o_2 _13078_ (.A1(\mem_state[0] ),
    .A2(mem_do_rinst),
    .B1(_10449_),
    .B2(_10447_),
    .C1(_10448_),
    .X(_10486_));
 sky130_fd_sc_hd__o311a_2 _13079_ (.A1(mem_do_wdata),
    .A2(_10484_),
    .A3(_10452_),
    .B1(_10485_),
    .C1(_10486_),
    .X(_10487_));
 sky130_fd_sc_hd__o21ai_2 _13080_ (.A1(_10482_),
    .A2(_10487_),
    .B1(_00300_),
    .Y(_10488_));
 sky130_vsdinv _13081_ (.A(_10488_),
    .Y(_10489_));
 sky130_fd_sc_hd__a32o_2 _13082_ (.A1(_12945_),
    .A2(_10480_),
    .A3(_10489_),
    .B1(\mem_state[1] ),
    .B2(_10488_),
    .X(_04068_));
 sky130_fd_sc_hd__a32o_2 _13083_ (.A1(_12944_),
    .A2(_10479_),
    .A3(_10489_),
    .B1(\mem_state[0] ),
    .B2(_10488_),
    .X(_04067_));
 sky130_vsdinv _13084_ (.A(mem_do_rinst),
    .Y(_10490_));
 sky130_fd_sc_hd__or2_2 _13085_ (.A(_10490_),
    .B(_10454_),
    .X(_10491_));
 sky130_vsdinv _13086_ (.A(_10491_),
    .Y(_10492_));
 sky130_fd_sc_hd__buf_1 _13087_ (.A(_10492_),
    .X(_10493_));
 sky130_fd_sc_hd__buf_1 _13088_ (.A(_10493_),
    .X(_12947_));
 sky130_fd_sc_hd__buf_1 _13089_ (.A(_10491_),
    .X(_10494_));
 sky130_fd_sc_hd__buf_1 _13090_ (.A(_10494_),
    .X(_00337_));
 sky130_vsdinv _13091_ (.A(_00327_),
    .Y(_10495_));
 sky130_fd_sc_hd__or3_2 _13092_ (.A(\mem_rdata_latched[28] ),
    .B(_10495_),
    .C(_00330_),
    .X(_10496_));
 sky130_vsdinv _13093_ (.A(_00325_),
    .Y(_10497_));
 sky130_vsdinv _13094_ (.A(_00324_),
    .Y(_10498_));
 sky130_fd_sc_hd__or3_2 _13095_ (.A(_10497_),
    .B(_10498_),
    .C(_00326_),
    .X(_10499_));
 sky130_fd_sc_hd__or4_2 _13096_ (.A(_00329_),
    .B(_00328_),
    .C(_10496_),
    .D(_10499_),
    .X(_10500_));
 sky130_fd_sc_hd__or2_2 _13097_ (.A(\mem_rdata_latched[27] ),
    .B(_10500_),
    .X(_10501_));
 sky130_fd_sc_hd__or3_2 _13098_ (.A(\mem_rdata_latched[31] ),
    .B(\mem_rdata_latched[30] ),
    .C(\mem_rdata_latched[29] ),
    .X(_10502_));
 sky130_fd_sc_hd__or3_2 _13099_ (.A(\mem_rdata_latched[26] ),
    .B(\mem_rdata_latched[25] ),
    .C(_10502_),
    .X(_10503_));
 sky130_fd_sc_hd__o21ba_2 _13100_ (.A1(_10501_),
    .A2(_10503_),
    .B1_N(\mem_rdata_latched[19] ),
    .X(_10504_));
 sky130_fd_sc_hd__or4b_2 _13101_ (.A(_10501_),
    .B(\mem_rdata_latched[25] ),
    .C(_10502_),
    .D_N(\mem_rdata_latched[26] ),
    .X(_10505_));
 sky130_vsdinv _13102_ (.A(\decoded_rs1[4] ),
    .Y(_00366_));
 sky130_fd_sc_hd__buf_1 _13103_ (.A(_10492_),
    .X(_10506_));
 sky130_fd_sc_hd__o22a_2 _13104_ (.A1(_10494_),
    .A2(_10505_),
    .B1(_00366_),
    .B2(_10506_),
    .X(_10507_));
 sky130_fd_sc_hd__o21ai_2 _13105_ (.A1(_00337_),
    .A2(_10504_),
    .B1(_10507_),
    .Y(_04066_));
 sky130_vsdinv _13106_ (.A(\cpu_state[1] ),
    .Y(_10508_));
 sky130_vsdinv _13107_ (.A(decoder_trigger),
    .Y(_10509_));
 sky130_vsdinv _13108_ (.A(\irq_mask[1] ),
    .Y(_10510_));
 sky130_vsdinv _13109_ (.A(\irq_mask[2] ),
    .Y(_10511_));
 sky130_vsdinv _13110_ (.A(\irq_pending[0] ),
    .Y(_10512_));
 sky130_vsdinv _13111_ (.A(\irq_pending[3] ),
    .Y(_10513_));
 sky130_fd_sc_hd__o22ai_2 _13112_ (.A1(\irq_mask[0] ),
    .A2(_10512_),
    .B1(\irq_mask[3] ),
    .B2(_10513_),
    .Y(_10514_));
 sky130_fd_sc_hd__a221o_2 _13113_ (.A1(_10510_),
    .A2(\irq_pending[1] ),
    .B1(_10511_),
    .B2(\irq_pending[2] ),
    .C1(_10514_),
    .X(_10515_));
 sky130_vsdinv _13114_ (.A(\irq_pending[17] ),
    .Y(_10516_));
 sky130_vsdinv _13115_ (.A(\irq_pending[19] ),
    .Y(_10517_));
 sky130_vsdinv _13116_ (.A(\irq_pending[16] ),
    .Y(_10518_));
 sky130_vsdinv _13117_ (.A(\irq_pending[18] ),
    .Y(_10519_));
 sky130_fd_sc_hd__o22a_2 _13118_ (.A1(\irq_mask[16] ),
    .A2(_10518_),
    .B1(\irq_mask[18] ),
    .B2(_10519_),
    .X(_10520_));
 sky130_fd_sc_hd__o221ai_2 _13119_ (.A1(\irq_mask[17] ),
    .A2(_10516_),
    .B1(\irq_mask[19] ),
    .B2(_10517_),
    .C1(_10520_),
    .Y(_10521_));
 sky130_vsdinv _13120_ (.A(\irq_mask[24] ),
    .Y(_10522_));
 sky130_vsdinv _13121_ (.A(\irq_mask[26] ),
    .Y(_10523_));
 sky130_vsdinv _13122_ (.A(\irq_pending[25] ),
    .Y(_10524_));
 sky130_vsdinv _13123_ (.A(\irq_pending[27] ),
    .Y(_10525_));
 sky130_fd_sc_hd__o22ai_2 _13124_ (.A1(\irq_mask[25] ),
    .A2(_10524_),
    .B1(\irq_mask[27] ),
    .B2(_10525_),
    .Y(_10526_));
 sky130_fd_sc_hd__a221o_2 _13125_ (.A1(_10522_),
    .A2(\irq_pending[24] ),
    .B1(_10523_),
    .B2(\irq_pending[26] ),
    .C1(_10526_),
    .X(_10527_));
 sky130_vsdinv _13126_ (.A(\irq_mask[5] ),
    .Y(_10528_));
 sky130_vsdinv _13127_ (.A(\irq_mask[7] ),
    .Y(_10529_));
 sky130_vsdinv _13128_ (.A(\irq_pending[4] ),
    .Y(_10530_));
 sky130_vsdinv _13129_ (.A(\irq_pending[6] ),
    .Y(_10531_));
 sky130_fd_sc_hd__o22ai_2 _13130_ (.A1(\irq_mask[4] ),
    .A2(_10530_),
    .B1(\irq_mask[6] ),
    .B2(_10531_),
    .Y(_10532_));
 sky130_fd_sc_hd__a221o_2 _13131_ (.A1(_10528_),
    .A2(\irq_pending[5] ),
    .B1(_10529_),
    .B2(\irq_pending[7] ),
    .C1(_10532_),
    .X(_10533_));
 sky130_fd_sc_hd__or4_4 _13132_ (.A(_10515_),
    .B(_10521_),
    .C(_10527_),
    .D(_10533_),
    .X(_10534_));
 sky130_vsdinv _13133_ (.A(\irq_mask[13] ),
    .Y(_10535_));
 sky130_vsdinv _13134_ (.A(\irq_mask[15] ),
    .Y(_10536_));
 sky130_vsdinv _13135_ (.A(\irq_pending[12] ),
    .Y(_10537_));
 sky130_vsdinv _13136_ (.A(\irq_pending[14] ),
    .Y(_10538_));
 sky130_fd_sc_hd__o22ai_2 _13137_ (.A1(\irq_mask[12] ),
    .A2(_10537_),
    .B1(\irq_mask[14] ),
    .B2(_10538_),
    .Y(_10539_));
 sky130_fd_sc_hd__a221o_2 _13138_ (.A1(_10535_),
    .A2(\irq_pending[13] ),
    .B1(_10536_),
    .B2(\irq_pending[15] ),
    .C1(_10539_),
    .X(_10540_));
 sky130_vsdinv _13139_ (.A(\irq_mask[28] ),
    .Y(_10541_));
 sky130_vsdinv _13140_ (.A(\irq_mask[30] ),
    .Y(_10542_));
 sky130_vsdinv _13141_ (.A(\irq_pending[29] ),
    .Y(_10543_));
 sky130_vsdinv _13142_ (.A(\irq_pending[31] ),
    .Y(_10544_));
 sky130_fd_sc_hd__o22ai_2 _13143_ (.A1(\irq_mask[29] ),
    .A2(_10543_),
    .B1(\irq_mask[31] ),
    .B2(_10544_),
    .Y(_10545_));
 sky130_fd_sc_hd__a221o_2 _13144_ (.A1(_10541_),
    .A2(\irq_pending[28] ),
    .B1(_10542_),
    .B2(\irq_pending[30] ),
    .C1(_10545_),
    .X(_10546_));
 sky130_vsdinv _13145_ (.A(\irq_mask[9] ),
    .Y(_10547_));
 sky130_vsdinv _13146_ (.A(\irq_mask[11] ),
    .Y(_10548_));
 sky130_vsdinv _13147_ (.A(\irq_pending[8] ),
    .Y(_10549_));
 sky130_vsdinv _13148_ (.A(\irq_pending[10] ),
    .Y(_10550_));
 sky130_fd_sc_hd__o22ai_2 _13149_ (.A1(\irq_mask[8] ),
    .A2(_10549_),
    .B1(\irq_mask[10] ),
    .B2(_10550_),
    .Y(_10551_));
 sky130_fd_sc_hd__a221o_2 _13150_ (.A1(_10547_),
    .A2(\irq_pending[9] ),
    .B1(_10548_),
    .B2(\irq_pending[11] ),
    .C1(_10551_),
    .X(_10552_));
 sky130_vsdinv _13151_ (.A(\irq_mask[20] ),
    .Y(_10553_));
 sky130_vsdinv _13152_ (.A(\irq_mask[22] ),
    .Y(_10554_));
 sky130_vsdinv _13153_ (.A(\irq_pending[21] ),
    .Y(_10555_));
 sky130_vsdinv _13154_ (.A(\irq_pending[23] ),
    .Y(_10556_));
 sky130_fd_sc_hd__o22ai_2 _13155_ (.A1(\irq_mask[21] ),
    .A2(_10555_),
    .B1(\irq_mask[23] ),
    .B2(_10556_),
    .Y(_10557_));
 sky130_fd_sc_hd__a221o_2 _13156_ (.A1(_10553_),
    .A2(\irq_pending[20] ),
    .B1(_10554_),
    .B2(\irq_pending[22] ),
    .C1(_10557_),
    .X(_10558_));
 sky130_fd_sc_hd__or4_4 _13157_ (.A(_10540_),
    .B(_10546_),
    .C(_10552_),
    .D(_10558_),
    .X(_10559_));
 sky130_vsdinv _13158_ (.A(irq_active),
    .Y(_10560_));
 sky130_vsdinv _13159_ (.A(irq_delay),
    .Y(_10561_));
 sky130_fd_sc_hd__o2111a_2 _13160_ (.A1(_10534_),
    .A2(_10559_),
    .B1(_10560_),
    .C1(_10561_),
    .D1(decoder_trigger),
    .X(_10562_));
 sky130_fd_sc_hd__or3_4 _13161_ (.A(\irq_state[1] ),
    .B(\irq_state[0] ),
    .C(_10562_),
    .X(_10563_));
 sky130_fd_sc_hd__o21ai_2 _13162_ (.A1(decoder_trigger),
    .A2(do_waitirq),
    .B1(instr_waitirq),
    .Y(_10564_));
 sky130_vsdinv _13163_ (.A(_10564_),
    .Y(_00309_));
 sky130_fd_sc_hd__or2_2 _13164_ (.A(_10563_),
    .B(_00309_),
    .X(_10565_));
 sky130_fd_sc_hd__or3_4 _13165_ (.A(_10508_),
    .B(_10509_),
    .C(_10565_),
    .X(_10566_));
 sky130_vsdinv _13166_ (.A(_10566_),
    .Y(_10567_));
 sky130_fd_sc_hd__o221a_2 _13167_ (.A1(irq_delay),
    .A2(_10567_),
    .B1(irq_active),
    .B2(_10566_),
    .C1(_10467_),
    .X(_04065_));
 sky130_vsdinv _13168_ (.A(pcpi_rs1[31]),
    .Y(_10568_));
 sky130_vsdinv _13169_ (.A(pcpi_valid),
    .Y(_10569_));
 sky130_fd_sc_hd__or2_2 _13170_ (.A(_10475_),
    .B(_10569_),
    .X(_10570_));
 sky130_fd_sc_hd__or4_2 _13171_ (.A(pcpi_insn[31]),
    .B(pcpi_insn[30]),
    .C(pcpi_insn[29]),
    .D(pcpi_insn[28]),
    .X(_10571_));
 sky130_fd_sc_hd__or4b_2 _13172_ (.A(pcpi_insn[27]),
    .B(pcpi_insn[26]),
    .C(pcpi_insn[14]),
    .D_N(pcpi_insn[25]),
    .X(_10572_));
 sky130_fd_sc_hd__or2b_2 _13173_ (.A(pcpi_insn[2]),
    .B_N(pcpi_insn[1]),
    .X(_10573_));
 sky130_fd_sc_hd__or4bb_2 _13174_ (.A(pcpi_insn[6]),
    .B(pcpi_insn[3]),
    .C_N(pcpi_insn[4]),
    .D_N(pcpi_insn[5]),
    .X(_10574_));
 sky130_fd_sc_hd__or4b_2 _13175_ (.A(_10572_),
    .B(_10573_),
    .C(_10574_),
    .D_N(pcpi_insn[0]),
    .X(_10575_));
 sky130_fd_sc_hd__or3_2 _13176_ (.A(_10570_),
    .B(_10571_),
    .C(_10575_),
    .X(_10576_));
 sky130_fd_sc_hd__or3_2 _13177_ (.A(\pcpi_mul.active[0] ),
    .B(\pcpi_mul.active[1] ),
    .C(_10576_),
    .X(_10577_));
 sky130_fd_sc_hd__buf_1 _13178_ (.A(_10577_),
    .X(_10578_));
 sky130_vsdinv _13179_ (.A(pcpi_insn[13]),
    .Y(_10579_));
 sky130_fd_sc_hd__or2b_2 _13180_ (.A(_10576_),
    .B_N(pcpi_insn[12]),
    .X(_10580_));
 sky130_vsdinv _13181_ (.A(_10580_),
    .Y(_10581_));
 sky130_fd_sc_hd__nor3_2 _13182_ (.A(_10579_),
    .B(pcpi_insn[12]),
    .C(_10576_),
    .Y(_10582_));
 sky130_fd_sc_hd__a21oi_2 _13183_ (.A1(_10579_),
    .A2(_10581_),
    .B1(_10582_),
    .Y(_10583_));
 sky130_vsdinv _13184_ (.A(\pcpi_mul.rs1[32] ),
    .Y(_10584_));
 sky130_fd_sc_hd__buf_1 _13185_ (.A(_10584_),
    .X(_10585_));
 sky130_fd_sc_hd__buf_1 _13186_ (.A(_10585_),
    .X(_10586_));
 sky130_fd_sc_hd__buf_1 _13187_ (.A(_10586_),
    .X(_10587_));
 sky130_fd_sc_hd__buf_1 _13188_ (.A(_10587_),
    .X(_10588_));
 sky130_fd_sc_hd__buf_1 _13189_ (.A(_10588_),
    .X(_10589_));
 sky130_vsdinv _13190_ (.A(_10577_),
    .Y(_10590_));
 sky130_fd_sc_hd__buf_1 _13191_ (.A(_10590_),
    .X(_10591_));
 sky130_fd_sc_hd__buf_1 _13192_ (.A(_10591_),
    .X(_10592_));
 sky130_fd_sc_hd__o32a_2 _13193_ (.A1(_10568_),
    .A2(_10578_),
    .A3(_10583_),
    .B1(_10589_),
    .B2(_10592_),
    .X(_10593_));
 sky130_vsdinv _13194_ (.A(_10593_),
    .Y(_04064_));
 sky130_vsdinv _13195_ (.A(pcpi_rs2[31]),
    .Y(_10594_));
 sky130_fd_sc_hd__or2_2 _13196_ (.A(pcpi_insn[13]),
    .B(_10580_),
    .X(_10595_));
 sky130_vsdinv _13197_ (.A(\pcpi_mul.rs2[32] ),
    .Y(_10596_));
 sky130_fd_sc_hd__buf_1 _13198_ (.A(_10596_),
    .X(_10597_));
 sky130_fd_sc_hd__buf_1 _13199_ (.A(_10597_),
    .X(_10598_));
 sky130_fd_sc_hd__buf_1 _13200_ (.A(_10598_),
    .X(_10599_));
 sky130_fd_sc_hd__buf_1 _13201_ (.A(_10599_),
    .X(_10600_));
 sky130_fd_sc_hd__buf_1 _13202_ (.A(_10590_),
    .X(_10601_));
 sky130_fd_sc_hd__o32a_2 _13203_ (.A1(_10594_),
    .A2(_10578_),
    .A3(_10595_),
    .B1(_10600_),
    .B2(_10601_),
    .X(_10602_));
 sky130_vsdinv _13204_ (.A(_10602_),
    .Y(_04063_));
 sky130_fd_sc_hd__buf_1 _13205_ (.A(\cpu_state[4] ),
    .X(_10603_));
 sky130_fd_sc_hd__buf_1 _13206_ (.A(_10603_),
    .X(_10604_));
 sky130_vsdinv _13207_ (.A(_00333_),
    .Y(_10605_));
 sky130_vsdinv _13208_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .Y(_10606_));
 sky130_fd_sc_hd__buf_1 _13209_ (.A(_10606_),
    .X(_10607_));
 sky130_fd_sc_hd__o21a_2 _13210_ (.A1(_10607_),
    .A2(alu_wait),
    .B1(_00333_),
    .X(_10608_));
 sky130_fd_sc_hd__o221a_2 _13211_ (.A1(_10604_),
    .A2(_10605_),
    .B1(latched_stalu),
    .B2(_10608_),
    .C1(_10467_),
    .X(_04062_));
 sky130_vsdinv _13212_ (.A(\cpu_state[4] ),
    .Y(_10609_));
 sky130_fd_sc_hd__buf_1 _13213_ (.A(_10609_),
    .X(_10610_));
 sky130_fd_sc_hd__inv_2 _13214_ (.A(alu_wait),
    .Y(_00302_));
 sky130_fd_sc_hd__or3_2 _13215_ (.A(\cpu_state[2] ),
    .B(\cpu_state[3] ),
    .C(\cpu_state[1] ),
    .X(_10611_));
 sky130_fd_sc_hd__or2_2 _13216_ (.A(_10603_),
    .B(_10457_),
    .X(_10612_));
 sky130_fd_sc_hd__or2_2 _13217_ (.A(_10611_),
    .B(_10612_),
    .X(_10613_));
 sky130_fd_sc_hd__buf_1 _13218_ (.A(\cpu_state[2] ),
    .X(_10614_));
 sky130_vsdinv _13219_ (.A(instr_rdcycle),
    .Y(_10615_));
 sky130_vsdinv _13220_ (.A(instr_rdinstrh),
    .Y(_10616_));
 sky130_vsdinv _13221_ (.A(instr_rdinstr),
    .Y(_10617_));
 sky130_vsdinv _13222_ (.A(instr_rdcycleh),
    .Y(_10618_));
 sky130_fd_sc_hd__and3_2 _13223_ (.A(_10616_),
    .B(_10617_),
    .C(_10618_),
    .X(_10619_));
 sky130_fd_sc_hd__buf_1 _13224_ (.A(_10619_),
    .X(_01714_));
 sky130_fd_sc_hd__or3_2 _13225_ (.A(instr_setq),
    .B(instr_getq),
    .C(instr_retirq),
    .X(_10620_));
 sky130_fd_sc_hd__nor3_2 _13226_ (.A(instr_maskirq),
    .B(_10620_),
    .C(instr_timer),
    .Y(_01717_));
 sky130_fd_sc_hd__and3_2 _13227_ (.A(_10615_),
    .B(_01714_),
    .C(_01717_),
    .X(_10621_));
 sky130_fd_sc_hd__nand2_2 _13228_ (.A(_10614_),
    .B(_10621_),
    .Y(_10622_));
 sky130_vsdinv _13229_ (.A(\pcpi_mul.active[1] ),
    .Y(_10623_));
 sky130_fd_sc_hd__nand2_2 _13230_ (.A(_10615_),
    .B(_01714_),
    .Y(_10624_));
 sky130_fd_sc_hd__or4_2 _13231_ (.A(instr_and),
    .B(instr_or),
    .C(instr_xor),
    .D(instr_sltu),
    .X(_10625_));
 sky130_fd_sc_hd__or4_2 _13232_ (.A(instr_sltiu),
    .B(instr_slti),
    .C(instr_bgeu),
    .D(instr_bge),
    .X(_10626_));
 sky130_fd_sc_hd__or4_2 _13233_ (.A(instr_maskirq),
    .B(_10620_),
    .C(_10625_),
    .D(_10626_),
    .X(_10627_));
 sky130_fd_sc_hd__or4_2 _13234_ (.A(instr_lw),
    .B(instr_lh),
    .C(instr_lb),
    .D(instr_jalr),
    .X(_10628_));
 sky130_fd_sc_hd__or4_2 _13235_ (.A(instr_sh),
    .B(instr_sb),
    .C(instr_lhu),
    .D(instr_lbu),
    .X(_10629_));
 sky130_fd_sc_hd__or2_2 _13236_ (.A(instr_auipc),
    .B(instr_lui),
    .X(_10630_));
 sky130_fd_sc_hd__or2_2 _13237_ (.A(instr_jal),
    .B(_10630_),
    .X(_00005_));
 sky130_fd_sc_hd__or4_2 _13238_ (.A(instr_sra),
    .B(instr_srai),
    .C(instr_srl),
    .D(instr_srli),
    .X(_10631_));
 sky130_fd_sc_hd__or4_2 _13239_ (.A(_10628_),
    .B(_10629_),
    .C(_00005_),
    .D(_10631_),
    .X(_10632_));
 sky130_fd_sc_hd__or4_2 _13240_ (.A(instr_andi),
    .B(instr_ori),
    .C(instr_xori),
    .D(instr_addi),
    .X(_10633_));
 sky130_fd_sc_hd__or4_2 _13241_ (.A(instr_slt),
    .B(instr_sll),
    .C(instr_sub),
    .D(instr_add),
    .X(_10634_));
 sky130_fd_sc_hd__or4_2 _13242_ (.A(instr_timer),
    .B(instr_waitirq),
    .C(instr_slli),
    .D(instr_sw),
    .X(_10635_));
 sky130_fd_sc_hd__or4_2 _13243_ (.A(instr_bltu),
    .B(instr_blt),
    .C(instr_bne),
    .D(instr_beq),
    .X(_10636_));
 sky130_fd_sc_hd__or4_2 _13244_ (.A(_10633_),
    .B(_10634_),
    .C(_10635_),
    .D(_10636_),
    .X(_10637_));
 sky130_fd_sc_hd__or4_2 _13245_ (.A(_10624_),
    .B(_10627_),
    .C(_10632_),
    .D(_10637_),
    .X(_10638_));
 sky130_fd_sc_hd__buf_1 _13246_ (.A(\cpu_state[3] ),
    .X(_10639_));
 sky130_fd_sc_hd__o21ai_2 _13247_ (.A1(_10623_),
    .A2(_10638_),
    .B1(_10639_),
    .Y(_10640_));
 sky130_fd_sc_hd__o2111a_2 _13248_ (.A1(_10610_),
    .A2(_00302_),
    .B1(_10613_),
    .C1(_10622_),
    .D1(_10640_),
    .X(_10641_));
 sky130_vsdinv _13249_ (.A(_10641_),
    .Y(_10642_));
 sky130_fd_sc_hd__o221a_2 _13250_ (.A1(_12981_),
    .A2(_10642_),
    .B1(latched_store),
    .B2(_10641_),
    .C1(_10467_),
    .X(_04061_));
 sky130_fd_sc_hd__buf_1 _13251_ (.A(_10482_),
    .X(_10643_));
 sky130_fd_sc_hd__buf_1 _13252_ (.A(_10643_),
    .X(_10644_));
 sky130_fd_sc_hd__buf_1 _13253_ (.A(\irq_state[1] ),
    .X(_10645_));
 sky130_fd_sc_hd__buf_1 _13254_ (.A(_10508_),
    .X(_10646_));
 sky130_fd_sc_hd__buf_1 _13255_ (.A(_10646_),
    .X(_10647_));
 sky130_vsdinv _13256_ (.A(\irq_state[0] ),
    .Y(_10648_));
 sky130_vsdinv _13257_ (.A(\irq_state[1] ),
    .Y(_10649_));
 sky130_fd_sc_hd__buf_1 _13258_ (.A(_10649_),
    .X(_10650_));
 sky130_fd_sc_hd__buf_1 _13259_ (.A(\cpu_state[1] ),
    .X(_10651_));
 sky130_fd_sc_hd__buf_1 _13260_ (.A(_10651_),
    .X(_10652_));
 sky130_fd_sc_hd__o32a_2 _13261_ (.A1(_10645_),
    .A2(_10647_),
    .A3(_10648_),
    .B1(_10650_),
    .B2(_10652_),
    .X(_10653_));
 sky130_fd_sc_hd__nor2_2 _13262_ (.A(_10644_),
    .B(_10653_),
    .Y(_04060_));
 sky130_fd_sc_hd__buf_1 _13263_ (.A(\irq_state[0] ),
    .X(_10654_));
 sky130_fd_sc_hd__buf_1 _13264_ (.A(_10654_),
    .X(_10655_));
 sky130_fd_sc_hd__buf_1 _13265_ (.A(_10655_),
    .X(_10656_));
 sky130_fd_sc_hd__buf_1 _13266_ (.A(_10652_),
    .X(_10657_));
 sky130_fd_sc_hd__buf_1 _13267_ (.A(_10463_),
    .X(_10658_));
 sky130_fd_sc_hd__a31o_2 _13268_ (.A1(_10649_),
    .A2(_10648_),
    .A3(_10562_),
    .B1(_10647_),
    .X(_10659_));
 sky130_fd_sc_hd__o211a_2 _13269_ (.A1(_10656_),
    .A2(_10657_),
    .B1(_10658_),
    .C1(_10659_),
    .X(_04059_));
 sky130_vsdinv _13270_ (.A(_00356_),
    .Y(_10660_));
 sky130_fd_sc_hd__or2_2 _13271_ (.A(_10475_),
    .B(_10453_),
    .X(_10661_));
 sky130_vsdinv _13272_ (.A(_10661_),
    .Y(_10662_));
 sky130_vsdinv _13273_ (.A(is_lb_lh_lw_lbu_lhu),
    .Y(_10663_));
 sky130_fd_sc_hd__inv_2 _13274_ (.A(_10638_),
    .Y(_00310_));
 sky130_fd_sc_hd__nor2_2 _13275_ (.A(_10663_),
    .B(_00310_),
    .Y(_10664_));
 sky130_fd_sc_hd__buf_1 _13276_ (.A(is_sb_sh_sw),
    .X(_10665_));
 sky130_vsdinv _13277_ (.A(_10665_),
    .Y(_10666_));
 sky130_fd_sc_hd__nor2_2 _13278_ (.A(_10666_),
    .B(_00310_),
    .Y(_10667_));
 sky130_fd_sc_hd__a22o_2 _13279_ (.A1(_10603_),
    .A2(alu_wait),
    .B1(_10609_),
    .B2(_10611_),
    .X(_10668_));
 sky130_fd_sc_hd__o221a_2 _13280_ (.A1(_10469_),
    .A2(_10664_),
    .B1(_10640_),
    .B2(_10667_),
    .C1(_10668_),
    .X(_10669_));
 sky130_fd_sc_hd__or2_2 _13281_ (.A(_10661_),
    .B(_10669_),
    .X(_10670_));
 sky130_fd_sc_hd__or2_2 _13282_ (.A(\cpu_state[6] ),
    .B(\cpu_state[5] ),
    .X(_10671_));
 sky130_fd_sc_hd__or4_2 _13283_ (.A(_10607_),
    .B(alu_wait),
    .C(_10481_),
    .D(_00343_),
    .X(_10672_));
 sky130_fd_sc_hd__nor4_2 _13284_ (.A(\cpu_state[0] ),
    .B(_10611_),
    .C(_10671_),
    .D(_10672_),
    .Y(_10673_));
 sky130_fd_sc_hd__nor2_2 _13285_ (.A(_10490_),
    .B(_10670_),
    .Y(_10674_));
 sky130_fd_sc_hd__a311o_2 _13286_ (.A1(_10660_),
    .A2(_10662_),
    .A3(_10670_),
    .B1(_10673_),
    .C1(_10674_),
    .X(_04058_));
 sky130_fd_sc_hd__or2_2 _13287_ (.A(instr_jal),
    .B(_10566_),
    .X(_10675_));
 sky130_vsdinv _13288_ (.A(_10675_),
    .Y(_10676_));
 sky130_fd_sc_hd__nor2_2 _13289_ (.A(instr_retirq),
    .B(instr_jalr),
    .Y(_10677_));
 sky130_fd_sc_hd__o221a_2 _13290_ (.A1(mem_do_prefetch),
    .A2(_10676_),
    .B1(_10675_),
    .B2(_10677_),
    .C1(_10662_),
    .X(_04057_));
 sky130_vsdinv _13291_ (.A(instr_maskirq),
    .Y(_10678_));
 sky130_fd_sc_hd__or2_2 _13292_ (.A(_10678_),
    .B(_10468_),
    .X(_10679_));
 sky130_fd_sc_hd__buf_1 _13293_ (.A(_10679_),
    .X(_10680_));
 sky130_fd_sc_hd__buf_1 _13294_ (.A(_10680_),
    .X(_10681_));
 sky130_fd_sc_hd__or3b_2 _13295_ (.A(_00362_),
    .B(_00360_),
    .C_N(_00368_),
    .X(_10682_));
 sky130_fd_sc_hd__or3_2 _13296_ (.A(_00358_),
    .B(_00357_),
    .C(_10682_),
    .X(_10683_));
 sky130_fd_sc_hd__inv_2 _13297_ (.A(_10683_),
    .Y(_10684_));
 sky130_fd_sc_hd__buf_1 _13298_ (.A(_10684_),
    .X(_10685_));
 sky130_fd_sc_hd__nor2_2 _13299_ (.A(_01207_),
    .B(_10685_),
    .Y(\cpuregs_rs1[31] ));
 sky130_vsdinv _13300_ (.A(_10679_),
    .Y(_10686_));
 sky130_fd_sc_hd__buf_1 _13301_ (.A(_10686_),
    .X(_10687_));
 sky130_fd_sc_hd__buf_1 _13302_ (.A(_10481_),
    .X(_10688_));
 sky130_fd_sc_hd__buf_1 _13303_ (.A(_10688_),
    .X(_10689_));
 sky130_fd_sc_hd__a221o_2 _13304_ (.A1(\irq_mask[31] ),
    .A2(_10681_),
    .B1(\cpuregs_rs1[31] ),
    .B2(_10687_),
    .C1(_10689_),
    .X(_04056_));
 sky130_fd_sc_hd__buf_1 _13305_ (.A(_10687_),
    .X(_10690_));
 sky130_fd_sc_hd__buf_1 _13306_ (.A(_10684_),
    .X(_10691_));
 sky130_fd_sc_hd__nor2_2 _13307_ (.A(_01180_),
    .B(_10691_),
    .Y(\cpuregs_rs1[30] ));
 sky130_fd_sc_hd__a221o_2 _13308_ (.A1(\irq_mask[30] ),
    .A2(_10681_),
    .B1(_10690_),
    .B2(\cpuregs_rs1[30] ),
    .C1(_10689_),
    .X(_04055_));
 sky130_fd_sc_hd__nor2_2 _13309_ (.A(_01153_),
    .B(_10685_),
    .Y(\cpuregs_rs1[29] ));
 sky130_fd_sc_hd__a221o_2 _13310_ (.A1(\irq_mask[29] ),
    .A2(_10681_),
    .B1(_10690_),
    .B2(\cpuregs_rs1[29] ),
    .C1(_10689_),
    .X(_04054_));
 sky130_fd_sc_hd__nor2_2 _13311_ (.A(_01126_),
    .B(_10691_),
    .Y(\cpuregs_rs1[28] ));
 sky130_fd_sc_hd__a221o_2 _13312_ (.A1(\irq_mask[28] ),
    .A2(_10681_),
    .B1(_10690_),
    .B2(\cpuregs_rs1[28] ),
    .C1(_10689_),
    .X(_04053_));
 sky130_fd_sc_hd__nor2_2 _13313_ (.A(_01099_),
    .B(_10685_),
    .Y(\cpuregs_rs1[27] ));
 sky130_fd_sc_hd__buf_1 _13314_ (.A(_10688_),
    .X(_10692_));
 sky130_fd_sc_hd__a221o_2 _13315_ (.A1(\irq_mask[27] ),
    .A2(_10681_),
    .B1(_10690_),
    .B2(\cpuregs_rs1[27] ),
    .C1(_10692_),
    .X(_04052_));
 sky130_fd_sc_hd__buf_1 _13316_ (.A(_10684_),
    .X(_10693_));
 sky130_fd_sc_hd__nor2_2 _13317_ (.A(_01072_),
    .B(_10693_),
    .Y(\cpuregs_rs1[26] ));
 sky130_fd_sc_hd__a221o_2 _13318_ (.A1(\irq_mask[26] ),
    .A2(_10681_),
    .B1(_10690_),
    .B2(\cpuregs_rs1[26] ),
    .C1(_10692_),
    .X(_04051_));
 sky130_fd_sc_hd__buf_1 _13319_ (.A(_10680_),
    .X(_10694_));
 sky130_fd_sc_hd__nor2_2 _13320_ (.A(_01045_),
    .B(_10685_),
    .Y(\cpuregs_rs1[25] ));
 sky130_fd_sc_hd__a221o_2 _13321_ (.A1(\irq_mask[25] ),
    .A2(_10694_),
    .B1(_10690_),
    .B2(\cpuregs_rs1[25] ),
    .C1(_10692_),
    .X(_04050_));
 sky130_fd_sc_hd__buf_1 _13322_ (.A(_10687_),
    .X(_10695_));
 sky130_fd_sc_hd__nor2_2 _13323_ (.A(_01018_),
    .B(_10693_),
    .Y(\cpuregs_rs1[24] ));
 sky130_fd_sc_hd__a221o_2 _13324_ (.A1(\irq_mask[24] ),
    .A2(_10694_),
    .B1(_10695_),
    .B2(\cpuregs_rs1[24] ),
    .C1(_10692_),
    .X(_04049_));
 sky130_fd_sc_hd__nor2_2 _13325_ (.A(_00991_),
    .B(_10685_),
    .Y(\cpuregs_rs1[23] ));
 sky130_fd_sc_hd__a221o_2 _13326_ (.A1(\irq_mask[23] ),
    .A2(_10694_),
    .B1(_10695_),
    .B2(\cpuregs_rs1[23] ),
    .C1(_10692_),
    .X(_04048_));
 sky130_fd_sc_hd__nor2_2 _13327_ (.A(_00964_),
    .B(_10693_),
    .Y(\cpuregs_rs1[22] ));
 sky130_fd_sc_hd__a221o_2 _13328_ (.A1(\irq_mask[22] ),
    .A2(_10694_),
    .B1(_10695_),
    .B2(\cpuregs_rs1[22] ),
    .C1(_10692_),
    .X(_04047_));
 sky130_fd_sc_hd__nor2_2 _13329_ (.A(_00937_),
    .B(_10685_),
    .Y(\cpuregs_rs1[21] ));
 sky130_fd_sc_hd__buf_1 _13330_ (.A(_10688_),
    .X(_10696_));
 sky130_fd_sc_hd__a221o_2 _13331_ (.A1(\irq_mask[21] ),
    .A2(_10694_),
    .B1(_10695_),
    .B2(\cpuregs_rs1[21] ),
    .C1(_10696_),
    .X(_04046_));
 sky130_fd_sc_hd__nor2_2 _13332_ (.A(_00910_),
    .B(_10693_),
    .Y(\cpuregs_rs1[20] ));
 sky130_fd_sc_hd__a221o_2 _13333_ (.A1(\irq_mask[20] ),
    .A2(_10694_),
    .B1(_10695_),
    .B2(\cpuregs_rs1[20] ),
    .C1(_10696_),
    .X(_04045_));
 sky130_fd_sc_hd__buf_1 _13334_ (.A(_10680_),
    .X(_10697_));
 sky130_fd_sc_hd__buf_1 _13335_ (.A(_10684_),
    .X(_10698_));
 sky130_fd_sc_hd__nor2_2 _13336_ (.A(_00883_),
    .B(_10698_),
    .Y(\cpuregs_rs1[19] ));
 sky130_fd_sc_hd__a221o_2 _13337_ (.A1(\irq_mask[19] ),
    .A2(_10697_),
    .B1(_10695_),
    .B2(\cpuregs_rs1[19] ),
    .C1(_10696_),
    .X(_04044_));
 sky130_fd_sc_hd__buf_1 _13338_ (.A(_10687_),
    .X(_10699_));
 sky130_fd_sc_hd__nor2_2 _13339_ (.A(_00856_),
    .B(_10693_),
    .Y(\cpuregs_rs1[18] ));
 sky130_fd_sc_hd__a221o_2 _13340_ (.A1(\irq_mask[18] ),
    .A2(_10697_),
    .B1(_10699_),
    .B2(\cpuregs_rs1[18] ),
    .C1(_10696_),
    .X(_04043_));
 sky130_fd_sc_hd__nor2_2 _13341_ (.A(_00829_),
    .B(_10698_),
    .Y(\cpuregs_rs1[17] ));
 sky130_fd_sc_hd__a221o_2 _13342_ (.A1(\irq_mask[17] ),
    .A2(_10697_),
    .B1(_10699_),
    .B2(\cpuregs_rs1[17] ),
    .C1(_10696_),
    .X(_04042_));
 sky130_fd_sc_hd__nor2_2 _13343_ (.A(_00802_),
    .B(_10698_),
    .Y(\cpuregs_rs1[16] ));
 sky130_fd_sc_hd__a221o_2 _13344_ (.A1(\irq_mask[16] ),
    .A2(_10697_),
    .B1(_10699_),
    .B2(\cpuregs_rs1[16] ),
    .C1(_10696_),
    .X(_04041_));
 sky130_fd_sc_hd__nor2_2 _13345_ (.A(_00775_),
    .B(_10693_),
    .Y(\cpuregs_rs1[15] ));
 sky130_fd_sc_hd__buf_1 _13346_ (.A(_10482_),
    .X(_10700_));
 sky130_fd_sc_hd__a221o_2 _13347_ (.A1(\irq_mask[15] ),
    .A2(_10697_),
    .B1(_10699_),
    .B2(\cpuregs_rs1[15] ),
    .C1(_10700_),
    .X(_04040_));
 sky130_fd_sc_hd__nor2_2 _13348_ (.A(_00748_),
    .B(_10698_),
    .Y(\cpuregs_rs1[14] ));
 sky130_fd_sc_hd__a221o_2 _13349_ (.A1(\irq_mask[14] ),
    .A2(_10697_),
    .B1(_10699_),
    .B2(\cpuregs_rs1[14] ),
    .C1(_10700_),
    .X(_04039_));
 sky130_fd_sc_hd__buf_1 _13350_ (.A(_10680_),
    .X(_10701_));
 sky130_fd_sc_hd__buf_1 _13351_ (.A(_10684_),
    .X(_10702_));
 sky130_fd_sc_hd__nor2_2 _13352_ (.A(_00721_),
    .B(_10702_),
    .Y(\cpuregs_rs1[13] ));
 sky130_fd_sc_hd__a221o_2 _13353_ (.A1(\irq_mask[13] ),
    .A2(_10701_),
    .B1(_10699_),
    .B2(\cpuregs_rs1[13] ),
    .C1(_10700_),
    .X(_04038_));
 sky130_fd_sc_hd__buf_1 _13354_ (.A(_10687_),
    .X(_10703_));
 sky130_fd_sc_hd__nor2_2 _13355_ (.A(_00694_),
    .B(_10698_),
    .Y(\cpuregs_rs1[12] ));
 sky130_fd_sc_hd__a221o_2 _13356_ (.A1(\irq_mask[12] ),
    .A2(_10701_),
    .B1(_10703_),
    .B2(\cpuregs_rs1[12] ),
    .C1(_10700_),
    .X(_04037_));
 sky130_fd_sc_hd__nor2_2 _13357_ (.A(_00667_),
    .B(_10702_),
    .Y(\cpuregs_rs1[11] ));
 sky130_fd_sc_hd__a221o_2 _13358_ (.A1(\irq_mask[11] ),
    .A2(_10701_),
    .B1(_10703_),
    .B2(\cpuregs_rs1[11] ),
    .C1(_10700_),
    .X(_04036_));
 sky130_fd_sc_hd__nor2_2 _13359_ (.A(_00640_),
    .B(_10698_),
    .Y(\cpuregs_rs1[10] ));
 sky130_fd_sc_hd__a221o_2 _13360_ (.A1(\irq_mask[10] ),
    .A2(_10701_),
    .B1(_10703_),
    .B2(\cpuregs_rs1[10] ),
    .C1(_10700_),
    .X(_04035_));
 sky130_fd_sc_hd__nor2_2 _13361_ (.A(_00613_),
    .B(_10702_),
    .Y(\cpuregs_rs1[9] ));
 sky130_fd_sc_hd__buf_1 _13362_ (.A(_10482_),
    .X(_10704_));
 sky130_fd_sc_hd__a221o_2 _13363_ (.A1(\irq_mask[9] ),
    .A2(_10701_),
    .B1(_10703_),
    .B2(\cpuregs_rs1[9] ),
    .C1(_10704_),
    .X(_04034_));
 sky130_fd_sc_hd__nor2_2 _13364_ (.A(_00586_),
    .B(_10691_),
    .Y(\cpuregs_rs1[8] ));
 sky130_fd_sc_hd__a221o_2 _13365_ (.A1(\irq_mask[8] ),
    .A2(_10701_),
    .B1(_10703_),
    .B2(\cpuregs_rs1[8] ),
    .C1(_10704_),
    .X(_04033_));
 sky130_fd_sc_hd__buf_1 _13366_ (.A(_10679_),
    .X(_10705_));
 sky130_fd_sc_hd__nor2_2 _13367_ (.A(_00559_),
    .B(_10702_),
    .Y(\cpuregs_rs1[7] ));
 sky130_fd_sc_hd__a221o_2 _13368_ (.A1(\irq_mask[7] ),
    .A2(_10705_),
    .B1(_10703_),
    .B2(\cpuregs_rs1[7] ),
    .C1(_10704_),
    .X(_04032_));
 sky130_fd_sc_hd__buf_1 _13369_ (.A(_10686_),
    .X(_10706_));
 sky130_fd_sc_hd__nor2_2 _13370_ (.A(_00532_),
    .B(_10691_),
    .Y(\cpuregs_rs1[6] ));
 sky130_fd_sc_hd__a221o_2 _13371_ (.A1(\irq_mask[6] ),
    .A2(_10705_),
    .B1(_10706_),
    .B2(\cpuregs_rs1[6] ),
    .C1(_10704_),
    .X(_04031_));
 sky130_fd_sc_hd__nor2_2 _13372_ (.A(_00505_),
    .B(_10702_),
    .Y(\cpuregs_rs1[5] ));
 sky130_fd_sc_hd__a221o_2 _13373_ (.A1(\irq_mask[5] ),
    .A2(_10705_),
    .B1(_10706_),
    .B2(\cpuregs_rs1[5] ),
    .C1(_10704_),
    .X(_04030_));
 sky130_fd_sc_hd__nor2_2 _13374_ (.A(_00478_),
    .B(_10691_),
    .Y(\cpuregs_rs1[4] ));
 sky130_fd_sc_hd__a221o_2 _13375_ (.A1(\irq_mask[4] ),
    .A2(_10705_),
    .B1(_10706_),
    .B2(\cpuregs_rs1[4] ),
    .C1(_10704_),
    .X(_04029_));
 sky130_fd_sc_hd__nor2_2 _13376_ (.A(_00451_),
    .B(_10691_),
    .Y(\cpuregs_rs1[3] ));
 sky130_fd_sc_hd__a221o_2 _13377_ (.A1(\irq_mask[3] ),
    .A2(_10705_),
    .B1(_10706_),
    .B2(\cpuregs_rs1[3] ),
    .C1(_10643_),
    .X(_04028_));
 sky130_fd_sc_hd__nor2_2 _13378_ (.A(_00424_),
    .B(_10702_),
    .Y(\cpuregs_rs1[2] ));
 sky130_fd_sc_hd__a221o_2 _13379_ (.A1(\irq_mask[2] ),
    .A2(_10705_),
    .B1(_10706_),
    .B2(\cpuregs_rs1[2] ),
    .C1(_10643_),
    .X(_04027_));
 sky130_fd_sc_hd__nor2_2 _13380_ (.A(_00397_),
    .B(_10684_),
    .Y(\cpuregs_rs1[1] ));
 sky130_fd_sc_hd__a221o_2 _13381_ (.A1(\irq_mask[1] ),
    .A2(_10680_),
    .B1(_10706_),
    .B2(\cpuregs_rs1[1] ),
    .C1(_10643_),
    .X(_04026_));
 sky130_fd_sc_hd__and2_2 _13382_ (.A(_00370_),
    .B(_10683_),
    .X(_10707_));
 sky130_fd_sc_hd__buf_1 _13383_ (.A(_10707_),
    .X(\cpuregs_rs1[0] ));
 sky130_fd_sc_hd__a221o_2 _13384_ (.A1(\irq_mask[0] ),
    .A2(_10680_),
    .B1(_10687_),
    .B2(\cpuregs_rs1[0] ),
    .C1(_10643_),
    .X(_04025_));
 sky130_vsdinv _13385_ (.A(mem_do_wdata),
    .Y(_10708_));
 sky130_fd_sc_hd__buf_1 _13386_ (.A(_10708_),
    .X(_00291_));
 sky130_fd_sc_hd__inv_2 _13387_ (.A(_10483_),
    .Y(_00301_));
 sky130_fd_sc_hd__a311o_2 _13388_ (.A1(_10456_),
    .A2(_00301_),
    .A3(_00291_),
    .B1(_10452_),
    .C1(_10476_),
    .X(_00316_));
 sky130_fd_sc_hd__or2_2 _13389_ (.A(trap),
    .B(_00316_),
    .X(_10709_));
 sky130_vsdinv _13390_ (.A(_10709_),
    .Y(_10710_));
 sky130_fd_sc_hd__buf_1 _13391_ (.A(_10709_),
    .X(_10711_));
 sky130_fd_sc_hd__buf_1 _13392_ (.A(_10711_),
    .X(_10712_));
 sky130_fd_sc_hd__a32o_2 _13393_ (.A1(_00291_),
    .A2(_10483_),
    .A3(_10710_),
    .B1(mem_instr),
    .B2(_10712_),
    .X(_04024_));
 sky130_vsdinv _13394_ (.A(_00329_),
    .Y(_10713_));
 sky130_fd_sc_hd__buf_1 _13395_ (.A(_00328_),
    .X(_10714_));
 sky130_fd_sc_hd__or3b_2 _13396_ (.A(_10713_),
    .B(_10714_),
    .C_N(_00330_),
    .X(_10715_));
 sky130_fd_sc_hd__nor3_2 _13397_ (.A(_00327_),
    .B(_10499_),
    .C(_10715_),
    .Y(_10716_));
 sky130_fd_sc_hd__o221a_2 _13398_ (.A1(_10494_),
    .A2(_10716_),
    .B1(is_beq_bne_blt_bge_bltu_bgeu),
    .B2(_10506_),
    .C1(_10467_),
    .X(_04023_));
 sky130_fd_sc_hd__buf_1 _13399_ (.A(_10492_),
    .X(_10717_));
 sky130_fd_sc_hd__buf_1 _13400_ (.A(_10491_),
    .X(_10718_));
 sky130_fd_sc_hd__buf_1 _13401_ (.A(_10718_),
    .X(_10719_));
 sky130_fd_sc_hd__a32o_2 _13402_ (.A1(\mem_rdata_latched[18] ),
    .A2(_10717_),
    .A3(_10505_),
    .B1(\decoded_rs1[3] ),
    .B2(_10719_),
    .X(_04022_));
 sky130_fd_sc_hd__a32o_2 _13403_ (.A1(\mem_rdata_latched[17] ),
    .A2(_10717_),
    .A3(_10505_),
    .B1(\decoded_rs1[2] ),
    .B2(_10719_),
    .X(_04021_));
 sky130_fd_sc_hd__a32o_2 _13404_ (.A1(\mem_rdata_latched[16] ),
    .A2(_10506_),
    .A3(_10505_),
    .B1(\decoded_rs1[1] ),
    .B2(_10719_),
    .X(_04020_));
 sky130_fd_sc_hd__a32o_2 _13405_ (.A1(\mem_rdata_latched[15] ),
    .A2(_10506_),
    .A3(_10505_),
    .B1(\decoded_rs1[0] ),
    .B2(_10719_),
    .X(_04019_));
 sky130_fd_sc_hd__or2_2 _13406_ (.A(_10509_),
    .B(decoder_pseudo_trigger),
    .X(_10720_));
 sky130_fd_sc_hd__buf_1 _13407_ (.A(_10720_),
    .X(_10721_));
 sky130_fd_sc_hd__buf_1 _13408_ (.A(_10721_),
    .X(_10722_));
 sky130_fd_sc_hd__buf_1 _13409_ (.A(_10722_),
    .X(_10723_));
 sky130_vsdinv _13410_ (.A(\mem_rdata_q[13] ),
    .Y(_10724_));
 sky130_fd_sc_hd__buf_1 _13411_ (.A(\mem_rdata_q[12] ),
    .X(_10725_));
 sky130_vsdinv _13412_ (.A(_10725_),
    .Y(_10726_));
 sky130_fd_sc_hd__buf_1 _13413_ (.A(\mem_rdata_q[14] ),
    .X(_10727_));
 sky130_vsdinv _13414_ (.A(_10727_),
    .Y(_10728_));
 sky130_fd_sc_hd__buf_1 _13415_ (.A(_10728_),
    .X(_00334_));
 sky130_fd_sc_hd__or3_2 _13416_ (.A(_10724_),
    .B(_10726_),
    .C(_00334_),
    .X(_10729_));
 sky130_vsdinv _13417_ (.A(is_alu_reg_reg),
    .Y(_10730_));
 sky130_fd_sc_hd__or4_2 _13418_ (.A(\mem_rdata_q[28] ),
    .B(\mem_rdata_q[26] ),
    .C(\mem_rdata_q[27] ),
    .D(\mem_rdata_q[25] ),
    .X(_10731_));
 sky130_fd_sc_hd__or4_2 _13419_ (.A(\mem_rdata_q[31] ),
    .B(\mem_rdata_q[30] ),
    .C(\mem_rdata_q[29] ),
    .D(_10731_),
    .X(_10732_));
 sky130_fd_sc_hd__or2_2 _13420_ (.A(_10720_),
    .B(_10732_),
    .X(_10733_));
 sky130_fd_sc_hd__or2_2 _13421_ (.A(_10730_),
    .B(_10733_),
    .X(_10734_));
 sky130_fd_sc_hd__o2bb2a_2 _13422_ (.A1_N(instr_and),
    .A2_N(_10723_),
    .B1(_10729_),
    .B2(_10734_),
    .X(_10735_));
 sky130_fd_sc_hd__nor2_2 _13423_ (.A(_10644_),
    .B(_10735_),
    .Y(_04018_));
 sky130_fd_sc_hd__or3_2 _13424_ (.A(_10724_),
    .B(_10725_),
    .C(_00334_),
    .X(_10736_));
 sky130_fd_sc_hd__o2bb2a_2 _13425_ (.A1_N(instr_or),
    .A2_N(_10723_),
    .B1(_10734_),
    .B2(_10736_),
    .X(_10737_));
 sky130_fd_sc_hd__nor2_2 _13426_ (.A(_10644_),
    .B(_10737_),
    .Y(_04017_));
 sky130_fd_sc_hd__buf_1 _13427_ (.A(\mem_rdata_q[13] ),
    .X(_10738_));
 sky130_fd_sc_hd__or3_2 _13428_ (.A(_10738_),
    .B(_10726_),
    .C(_10728_),
    .X(_10739_));
 sky130_fd_sc_hd__buf_1 _13429_ (.A(\mem_rdata_q[29] ),
    .X(_10740_));
 sky130_fd_sc_hd__buf_1 _13430_ (.A(_10721_),
    .X(_10741_));
 sky130_fd_sc_hd__buf_1 _13431_ (.A(\mem_rdata_q[31] ),
    .X(_10742_));
 sky130_vsdinv _13432_ (.A(\mem_rdata_q[30] ),
    .Y(_10743_));
 sky130_fd_sc_hd__or3_2 _13433_ (.A(_10742_),
    .B(_10743_),
    .C(_10731_),
    .X(_10744_));
 sky130_fd_sc_hd__or3_2 _13434_ (.A(_10740_),
    .B(_10741_),
    .C(_10744_),
    .X(_10745_));
 sky130_vsdinv _13435_ (.A(instr_sra),
    .Y(_10746_));
 sky130_vsdinv _13436_ (.A(_10721_),
    .Y(_10747_));
 sky130_fd_sc_hd__buf_1 _13437_ (.A(_10747_),
    .X(_10748_));
 sky130_fd_sc_hd__buf_1 _13438_ (.A(_10748_),
    .X(_10749_));
 sky130_fd_sc_hd__o32a_2 _13439_ (.A1(_10730_),
    .A2(_10739_),
    .A3(_10745_),
    .B1(_10746_),
    .B2(_10749_),
    .X(_10750_));
 sky130_fd_sc_hd__nor2_2 _13440_ (.A(_10644_),
    .B(_10750_),
    .Y(_04016_));
 sky130_vsdinv _13441_ (.A(instr_srl),
    .Y(_10751_));
 sky130_fd_sc_hd__o32a_2 _13442_ (.A1(_10730_),
    .A2(_10739_),
    .A3(_10733_),
    .B1(_10751_),
    .B2(_10749_),
    .X(_10752_));
 sky130_fd_sc_hd__nor2_2 _13443_ (.A(_10644_),
    .B(_10752_),
    .Y(_04015_));
 sky130_fd_sc_hd__or3_2 _13444_ (.A(_10738_),
    .B(_10725_),
    .C(_00334_),
    .X(_10753_));
 sky130_fd_sc_hd__o2bb2a_2 _13445_ (.A1_N(instr_xor),
    .A2_N(_10723_),
    .B1(_10734_),
    .B2(_10753_),
    .X(_10754_));
 sky130_fd_sc_hd__nor2_2 _13446_ (.A(_10644_),
    .B(_10754_),
    .Y(_04014_));
 sky130_fd_sc_hd__buf_1 _13447_ (.A(_10643_),
    .X(_10755_));
 sky130_fd_sc_hd__or3_2 _13448_ (.A(_10724_),
    .B(_10726_),
    .C(_10727_),
    .X(_10756_));
 sky130_fd_sc_hd__o2bb2a_2 _13449_ (.A1_N(instr_sltu),
    .A2_N(_10723_),
    .B1(_10734_),
    .B2(_10756_),
    .X(_10757_));
 sky130_fd_sc_hd__nor2_2 _13450_ (.A(_10755_),
    .B(_10757_),
    .Y(_04013_));
 sky130_fd_sc_hd__or3_2 _13451_ (.A(_10724_),
    .B(\mem_rdata_q[12] ),
    .C(\mem_rdata_q[14] ),
    .X(_10758_));
 sky130_fd_sc_hd__o2bb2a_2 _13452_ (.A1_N(instr_slt),
    .A2_N(_10723_),
    .B1(_10734_),
    .B2(_10758_),
    .X(_10759_));
 sky130_fd_sc_hd__nor2_2 _13453_ (.A(_10755_),
    .B(_10759_),
    .Y(_04012_));
 sky130_fd_sc_hd__buf_1 _13454_ (.A(_10741_),
    .X(_10760_));
 sky130_fd_sc_hd__or3_2 _13455_ (.A(_10738_),
    .B(_10726_),
    .C(_10727_),
    .X(_10761_));
 sky130_fd_sc_hd__o2bb2a_2 _13456_ (.A1_N(instr_sll),
    .A2_N(_10760_),
    .B1(_10734_),
    .B2(_10761_),
    .X(_10762_));
 sky130_fd_sc_hd__nor2_2 _13457_ (.A(_10755_),
    .B(_10762_),
    .Y(_04011_));
 sky130_fd_sc_hd__or3_2 _13458_ (.A(\mem_rdata_q[13] ),
    .B(_10725_),
    .C(_10727_),
    .X(_10763_));
 sky130_vsdinv _13459_ (.A(instr_sub),
    .Y(_10764_));
 sky130_fd_sc_hd__o32a_2 _13460_ (.A1(_10730_),
    .A2(_10763_),
    .A3(_10745_),
    .B1(_10764_),
    .B2(_10749_),
    .X(_10765_));
 sky130_fd_sc_hd__nor2_2 _13461_ (.A(_10755_),
    .B(_10765_),
    .Y(_04010_));
 sky130_vsdinv _13462_ (.A(instr_add),
    .Y(_10766_));
 sky130_fd_sc_hd__o32a_2 _13463_ (.A1(_10730_),
    .A2(_10763_),
    .A3(_10733_),
    .B1(_10766_),
    .B2(_10749_),
    .X(_10767_));
 sky130_fd_sc_hd__nor2_2 _13464_ (.A(_10755_),
    .B(_10767_),
    .Y(_04009_));
 sky130_vsdinv _13465_ (.A(is_alu_reg_imm),
    .Y(_10768_));
 sky130_fd_sc_hd__buf_1 _13466_ (.A(_10768_),
    .X(_10769_));
 sky130_fd_sc_hd__buf_1 _13467_ (.A(_10741_),
    .X(_10770_));
 sky130_vsdinv _13468_ (.A(instr_andi),
    .Y(_10771_));
 sky130_fd_sc_hd__buf_1 _13469_ (.A(_10748_),
    .X(_10772_));
 sky130_fd_sc_hd__o32a_2 _13470_ (.A1(_10769_),
    .A2(_10770_),
    .A3(_10729_),
    .B1(_10771_),
    .B2(_10772_),
    .X(_10773_));
 sky130_fd_sc_hd__nor2_2 _13471_ (.A(_10755_),
    .B(_10773_),
    .Y(_04008_));
 sky130_fd_sc_hd__buf_1 _13472_ (.A(_10481_),
    .X(_10774_));
 sky130_fd_sc_hd__buf_1 _13473_ (.A(_10774_),
    .X(_10775_));
 sky130_vsdinv _13474_ (.A(instr_ori),
    .Y(_10776_));
 sky130_fd_sc_hd__o32a_2 _13475_ (.A1(_10769_),
    .A2(_10770_),
    .A3(_10736_),
    .B1(_10776_),
    .B2(_10772_),
    .X(_10777_));
 sky130_fd_sc_hd__nor2_2 _13476_ (.A(_10775_),
    .B(_10777_),
    .Y(_04007_));
 sky130_vsdinv _13477_ (.A(instr_xori),
    .Y(_10778_));
 sky130_fd_sc_hd__o32a_2 _13478_ (.A1(_10769_),
    .A2(_10770_),
    .A3(_10753_),
    .B1(_10778_),
    .B2(_10772_),
    .X(_10779_));
 sky130_fd_sc_hd__nor2_2 _13479_ (.A(_10775_),
    .B(_10779_),
    .Y(_04006_));
 sky130_vsdinv _13480_ (.A(instr_sltiu),
    .Y(_10780_));
 sky130_fd_sc_hd__o32a_2 _13481_ (.A1(_10769_),
    .A2(_10770_),
    .A3(_10756_),
    .B1(_10780_),
    .B2(_10772_),
    .X(_10781_));
 sky130_fd_sc_hd__nor2_2 _13482_ (.A(_10775_),
    .B(_10781_),
    .Y(_04005_));
 sky130_vsdinv _13483_ (.A(instr_slti),
    .Y(_10782_));
 sky130_fd_sc_hd__o32a_2 _13484_ (.A1(_10768_),
    .A2(_10770_),
    .A3(_10758_),
    .B1(_10782_),
    .B2(_10772_),
    .X(_10783_));
 sky130_fd_sc_hd__nor2_2 _13485_ (.A(_10775_),
    .B(_10783_),
    .Y(_04004_));
 sky130_vsdinv _13486_ (.A(instr_addi),
    .Y(_10784_));
 sky130_fd_sc_hd__o32a_2 _13487_ (.A1(_10768_),
    .A2(_10770_),
    .A3(_10763_),
    .B1(_10784_),
    .B2(_10772_),
    .X(_10785_));
 sky130_fd_sc_hd__nor2_2 _13488_ (.A(_10775_),
    .B(_10785_),
    .Y(_04003_));
 sky130_fd_sc_hd__buf_1 _13489_ (.A(_10607_),
    .X(_10786_));
 sky130_fd_sc_hd__buf_1 _13490_ (.A(_10741_),
    .X(_10787_));
 sky130_vsdinv _13491_ (.A(instr_bgeu),
    .Y(_10788_));
 sky130_fd_sc_hd__buf_1 _13492_ (.A(_10748_),
    .X(_10789_));
 sky130_fd_sc_hd__o32a_2 _13493_ (.A1(_10786_),
    .A2(_10787_),
    .A3(_10729_),
    .B1(_10788_),
    .B2(_10789_),
    .X(_10790_));
 sky130_fd_sc_hd__nor2_2 _13494_ (.A(_10775_),
    .B(_10790_),
    .Y(_04002_));
 sky130_fd_sc_hd__buf_1 _13495_ (.A(_10774_),
    .X(_10791_));
 sky130_vsdinv _13496_ (.A(instr_bltu),
    .Y(_10792_));
 sky130_fd_sc_hd__o32a_2 _13497_ (.A1(_10786_),
    .A2(_10787_),
    .A3(_10736_),
    .B1(_10792_),
    .B2(_10789_),
    .X(_10793_));
 sky130_fd_sc_hd__nor2_2 _13498_ (.A(_10791_),
    .B(_10793_),
    .Y(_04001_));
 sky130_vsdinv _13499_ (.A(instr_bge),
    .Y(_10794_));
 sky130_fd_sc_hd__o32a_2 _13500_ (.A1(_10786_),
    .A2(_10787_),
    .A3(_10739_),
    .B1(_10794_),
    .B2(_10789_),
    .X(_10795_));
 sky130_fd_sc_hd__nor2_2 _13501_ (.A(_10791_),
    .B(_10795_),
    .Y(_04000_));
 sky130_vsdinv _13502_ (.A(instr_blt),
    .Y(_10796_));
 sky130_fd_sc_hd__o32a_2 _13503_ (.A1(_10786_),
    .A2(_10787_),
    .A3(_10753_),
    .B1(_10796_),
    .B2(_10789_),
    .X(_10797_));
 sky130_fd_sc_hd__nor2_2 _13504_ (.A(_10791_),
    .B(_10797_),
    .Y(_03999_));
 sky130_vsdinv _13505_ (.A(instr_bne),
    .Y(_10798_));
 sky130_fd_sc_hd__o32a_2 _13506_ (.A1(_10786_),
    .A2(_10787_),
    .A3(_10761_),
    .B1(_10798_),
    .B2(_10789_),
    .X(_10799_));
 sky130_fd_sc_hd__nor2_2 _13507_ (.A(_10791_),
    .B(_10799_),
    .Y(_03998_));
 sky130_vsdinv _13508_ (.A(instr_beq),
    .Y(_10800_));
 sky130_fd_sc_hd__o32a_2 _13509_ (.A1(_10607_),
    .A2(_10787_),
    .A3(_10763_),
    .B1(_10800_),
    .B2(_10789_),
    .X(_10801_));
 sky130_fd_sc_hd__nor2_2 _13510_ (.A(_10791_),
    .B(_10801_),
    .Y(_03997_));
 sky130_fd_sc_hd__or2_2 _13511_ (.A(\pcpi_timeout_counter[1] ),
    .B(\pcpi_timeout_counter[0] ),
    .X(_10802_));
 sky130_fd_sc_hd__or2_2 _13512_ (.A(\pcpi_timeout_counter[2] ),
    .B(_10802_),
    .X(_10803_));
 sky130_fd_sc_hd__a21o_2 _13513_ (.A1(\pcpi_timeout_counter[3] ),
    .A2(_10803_),
    .B1(_10570_),
    .X(_03996_));
 sky130_vsdinv _13514_ (.A(_10803_),
    .Y(_10804_));
 sky130_fd_sc_hd__a221o_2 _13515_ (.A1(\pcpi_timeout_counter[2] ),
    .A2(_10802_),
    .B1(\pcpi_timeout_counter[3] ),
    .B2(_10804_),
    .C1(_10570_),
    .X(_03995_));
 sky130_vsdinv _13516_ (.A(_10802_),
    .Y(_10805_));
 sky130_fd_sc_hd__or2_2 _13517_ (.A(\pcpi_timeout_counter[3] ),
    .B(_10803_),
    .X(_10806_));
 sky130_fd_sc_hd__a221o_2 _13518_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(\pcpi_timeout_counter[0] ),
    .B1(_10805_),
    .B2(_10806_),
    .C1(_10570_),
    .X(_03994_));
 sky130_vsdinv _13519_ (.A(\pcpi_timeout_counter[0] ),
    .Y(_10807_));
 sky130_fd_sc_hd__a21o_2 _13520_ (.A1(_10807_),
    .A2(_10806_),
    .B1(_10570_),
    .X(_03993_));
 sky130_vsdinv _13521_ (.A(_10455_),
    .Y(_10808_));
 sky130_fd_sc_hd__buf_1 _13522_ (.A(_10808_),
    .X(_00296_));
 sky130_fd_sc_hd__or2_2 _13523_ (.A(_10476_),
    .B(mem_do_wdata),
    .X(_10809_));
 sky130_fd_sc_hd__or4_2 _13524_ (.A(\cpu_state[0] ),
    .B(_10611_),
    .C(_10612_),
    .D(_10809_),
    .X(_10810_));
 sky130_fd_sc_hd__o22ai_2 _13525_ (.A1(_00291_),
    .A2(_10661_),
    .B1(_00296_),
    .B2(_10810_),
    .Y(_03992_));
 sky130_fd_sc_hd__buf_1 _13526_ (.A(_10456_),
    .X(_10811_));
 sky130_fd_sc_hd__or3_2 _13527_ (.A(_10477_),
    .B(mem_do_rdata),
    .C(_10458_),
    .X(_10812_));
 sky130_fd_sc_hd__o22ai_2 _13528_ (.A1(_10811_),
    .A2(_10661_),
    .B1(_00296_),
    .B2(_10812_),
    .Y(_03991_));
 sky130_fd_sc_hd__buf_1 _13529_ (.A(_10646_),
    .X(_10813_));
 sky130_fd_sc_hd__buf_1 _13530_ (.A(_10466_),
    .X(_10814_));
 sky130_fd_sc_hd__o221a_2 _13531_ (.A1(\reg_next_pc[31] ),
    .A2(_10652_),
    .B1(_02530_),
    .B2(_10813_),
    .C1(_10814_),
    .X(_03990_));
 sky130_fd_sc_hd__buf_1 _13532_ (.A(_10647_),
    .X(_00322_));
 sky130_fd_sc_hd__o221a_2 _13533_ (.A1(_10657_),
    .A2(\reg_next_pc[30] ),
    .B1(_00322_),
    .B2(_02529_),
    .C1(_10814_),
    .X(_03989_));
 sky130_fd_sc_hd__o221a_2 _13534_ (.A1(_10657_),
    .A2(\reg_next_pc[29] ),
    .B1(_00322_),
    .B2(_02527_),
    .C1(_10814_),
    .X(_03988_));
 sky130_fd_sc_hd__buf_1 _13535_ (.A(_10647_),
    .X(_10815_));
 sky130_fd_sc_hd__o221a_2 _13536_ (.A1(_10657_),
    .A2(\reg_next_pc[28] ),
    .B1(_10815_),
    .B2(_02526_),
    .C1(_10814_),
    .X(_03987_));
 sky130_fd_sc_hd__o221a_2 _13537_ (.A1(_10657_),
    .A2(\reg_next_pc[27] ),
    .B1(_10815_),
    .B2(_02525_),
    .C1(_10814_),
    .X(_03986_));
 sky130_fd_sc_hd__o221a_2 _13538_ (.A1(_10657_),
    .A2(\reg_next_pc[26] ),
    .B1(_10815_),
    .B2(_02524_),
    .C1(_10814_),
    .X(_03985_));
 sky130_fd_sc_hd__buf_1 _13539_ (.A(_10651_),
    .X(_10816_));
 sky130_fd_sc_hd__buf_1 _13540_ (.A(_10816_),
    .X(_10817_));
 sky130_fd_sc_hd__buf_1 _13541_ (.A(_10466_),
    .X(_10818_));
 sky130_fd_sc_hd__o221a_2 _13542_ (.A1(_10817_),
    .A2(\reg_next_pc[25] ),
    .B1(_10815_),
    .B2(_02523_),
    .C1(_10818_),
    .X(_03984_));
 sky130_fd_sc_hd__o221a_2 _13543_ (.A1(_10817_),
    .A2(\reg_next_pc[24] ),
    .B1(_10815_),
    .B2(_02522_),
    .C1(_10818_),
    .X(_03983_));
 sky130_fd_sc_hd__o221a_2 _13544_ (.A1(_10817_),
    .A2(\reg_next_pc[23] ),
    .B1(_10815_),
    .B2(_02521_),
    .C1(_10818_),
    .X(_03982_));
 sky130_fd_sc_hd__buf_1 _13545_ (.A(_10647_),
    .X(_10819_));
 sky130_fd_sc_hd__o221a_2 _13546_ (.A1(_10817_),
    .A2(\reg_next_pc[22] ),
    .B1(_10819_),
    .B2(_02520_),
    .C1(_10818_),
    .X(_03981_));
 sky130_fd_sc_hd__o221a_2 _13547_ (.A1(_10817_),
    .A2(\reg_next_pc[21] ),
    .B1(_10819_),
    .B2(_02519_),
    .C1(_10818_),
    .X(_03980_));
 sky130_fd_sc_hd__o221a_2 _13548_ (.A1(_10817_),
    .A2(\reg_next_pc[20] ),
    .B1(_10819_),
    .B2(_02518_),
    .C1(_10818_),
    .X(_03979_));
 sky130_fd_sc_hd__buf_1 _13549_ (.A(_10816_),
    .X(_10820_));
 sky130_fd_sc_hd__buf_1 _13550_ (.A(_10466_),
    .X(_10821_));
 sky130_fd_sc_hd__o221a_2 _13551_ (.A1(_10820_),
    .A2(\reg_next_pc[19] ),
    .B1(_10819_),
    .B2(_02516_),
    .C1(_10821_),
    .X(_03978_));
 sky130_fd_sc_hd__o221a_2 _13552_ (.A1(_10820_),
    .A2(\reg_next_pc[18] ),
    .B1(_10819_),
    .B2(_02515_),
    .C1(_10821_),
    .X(_03977_));
 sky130_fd_sc_hd__o221a_2 _13553_ (.A1(_10820_),
    .A2(\reg_next_pc[17] ),
    .B1(_10819_),
    .B2(_02514_),
    .C1(_10821_),
    .X(_03976_));
 sky130_fd_sc_hd__buf_1 _13554_ (.A(_10647_),
    .X(_10822_));
 sky130_fd_sc_hd__o221a_2 _13555_ (.A1(_10820_),
    .A2(\reg_next_pc[16] ),
    .B1(_10822_),
    .B2(_02513_),
    .C1(_10821_),
    .X(_03975_));
 sky130_fd_sc_hd__o221a_2 _13556_ (.A1(_10820_),
    .A2(\reg_next_pc[15] ),
    .B1(_10822_),
    .B2(_02512_),
    .C1(_10821_),
    .X(_03974_));
 sky130_fd_sc_hd__o221a_2 _13557_ (.A1(_10820_),
    .A2(\reg_next_pc[14] ),
    .B1(_10822_),
    .B2(_02511_),
    .C1(_10821_),
    .X(_03973_));
 sky130_fd_sc_hd__buf_1 _13558_ (.A(_10816_),
    .X(_10823_));
 sky130_fd_sc_hd__buf_1 _13559_ (.A(_10466_),
    .X(_10824_));
 sky130_fd_sc_hd__o221a_2 _13560_ (.A1(_10823_),
    .A2(\reg_next_pc[13] ),
    .B1(_10822_),
    .B2(_02510_),
    .C1(_10824_),
    .X(_03972_));
 sky130_fd_sc_hd__o221a_2 _13561_ (.A1(_10823_),
    .A2(\reg_next_pc[12] ),
    .B1(_10822_),
    .B2(_02509_),
    .C1(_10824_),
    .X(_03971_));
 sky130_fd_sc_hd__o221a_2 _13562_ (.A1(_10823_),
    .A2(\reg_next_pc[11] ),
    .B1(_10822_),
    .B2(_02508_),
    .C1(_10824_),
    .X(_03970_));
 sky130_fd_sc_hd__buf_1 _13563_ (.A(_10646_),
    .X(_10825_));
 sky130_fd_sc_hd__buf_1 _13564_ (.A(_10825_),
    .X(_10826_));
 sky130_fd_sc_hd__o221a_2 _13565_ (.A1(_10823_),
    .A2(\reg_next_pc[10] ),
    .B1(_10826_),
    .B2(_02507_),
    .C1(_10824_),
    .X(_03969_));
 sky130_fd_sc_hd__o221a_2 _13566_ (.A1(_10823_),
    .A2(\reg_next_pc[9] ),
    .B1(_10826_),
    .B2(_02537_),
    .C1(_10824_),
    .X(_03968_));
 sky130_fd_sc_hd__o221a_2 _13567_ (.A1(_10823_),
    .A2(\reg_next_pc[8] ),
    .B1(_10826_),
    .B2(_02536_),
    .C1(_10824_),
    .X(_03967_));
 sky130_fd_sc_hd__buf_1 _13568_ (.A(_10816_),
    .X(_10827_));
 sky130_fd_sc_hd__buf_1 _13569_ (.A(_10444_),
    .X(_10828_));
 sky130_fd_sc_hd__buf_1 _13570_ (.A(_10828_),
    .X(_10829_));
 sky130_fd_sc_hd__o221a_2 _13571_ (.A1(_10827_),
    .A2(\reg_next_pc[7] ),
    .B1(_10826_),
    .B2(_02535_),
    .C1(_10829_),
    .X(_03966_));
 sky130_fd_sc_hd__o221a_2 _13572_ (.A1(_10827_),
    .A2(\reg_next_pc[6] ),
    .B1(_10826_),
    .B2(_02534_),
    .C1(_10829_),
    .X(_03965_));
 sky130_fd_sc_hd__o221a_2 _13573_ (.A1(_10827_),
    .A2(\reg_next_pc[5] ),
    .B1(_10826_),
    .B2(_02533_),
    .C1(_10829_),
    .X(_03964_));
 sky130_fd_sc_hd__buf_1 _13574_ (.A(_10825_),
    .X(_10830_));
 sky130_fd_sc_hd__o221a_2 _13575_ (.A1(_10827_),
    .A2(\reg_next_pc[4] ),
    .B1(_10830_),
    .B2(_02532_),
    .C1(_10829_),
    .X(_03963_));
 sky130_fd_sc_hd__o221a_2 _13576_ (.A1(_10827_),
    .A2(\reg_next_pc[3] ),
    .B1(_10830_),
    .B2(_02531_),
    .C1(_10829_),
    .X(_03962_));
 sky130_fd_sc_hd__o221a_2 _13577_ (.A1(_10827_),
    .A2(\reg_next_pc[2] ),
    .B1(_10830_),
    .B2(_02528_),
    .C1(_10829_),
    .X(_03961_));
 sky130_fd_sc_hd__buf_1 _13578_ (.A(_10816_),
    .X(_10831_));
 sky130_fd_sc_hd__buf_1 _13579_ (.A(_10828_),
    .X(_10832_));
 sky130_fd_sc_hd__o221a_2 _13580_ (.A1(_10831_),
    .A2(\reg_next_pc[1] ),
    .B1(_10830_),
    .B2(_02517_),
    .C1(_10832_),
    .X(_03960_));
 sky130_fd_sc_hd__o221a_2 _13581_ (.A1(_10831_),
    .A2(\reg_pc[31] ),
    .B1(_10830_),
    .B2(_02581_),
    .C1(_10832_),
    .X(_03959_));
 sky130_fd_sc_hd__o221a_2 _13582_ (.A1(_10831_),
    .A2(\reg_pc[30] ),
    .B1(_10830_),
    .B2(_02580_),
    .C1(_10832_),
    .X(_03958_));
 sky130_fd_sc_hd__buf_1 _13583_ (.A(_10825_),
    .X(_10833_));
 sky130_fd_sc_hd__o221a_2 _13584_ (.A1(_10831_),
    .A2(\reg_pc[29] ),
    .B1(_10833_),
    .B2(_02579_),
    .C1(_10832_),
    .X(_03957_));
 sky130_fd_sc_hd__o221a_2 _13585_ (.A1(_10831_),
    .A2(\reg_pc[28] ),
    .B1(_10833_),
    .B2(_02578_),
    .C1(_10832_),
    .X(_03956_));
 sky130_fd_sc_hd__o221a_2 _13586_ (.A1(_10831_),
    .A2(\reg_pc[27] ),
    .B1(_10833_),
    .B2(_02577_),
    .C1(_10832_),
    .X(_03955_));
 sky130_fd_sc_hd__buf_1 _13587_ (.A(_10816_),
    .X(_10834_));
 sky130_fd_sc_hd__buf_1 _13588_ (.A(_10828_),
    .X(_10835_));
 sky130_fd_sc_hd__o221a_2 _13589_ (.A1(_10834_),
    .A2(\reg_pc[26] ),
    .B1(_10833_),
    .B2(_02576_),
    .C1(_10835_),
    .X(_03954_));
 sky130_fd_sc_hd__o221a_2 _13590_ (.A1(_10834_),
    .A2(\reg_pc[25] ),
    .B1(_10833_),
    .B2(_02575_),
    .C1(_10835_),
    .X(_03953_));
 sky130_fd_sc_hd__o221a_2 _13591_ (.A1(_10834_),
    .A2(\reg_pc[24] ),
    .B1(_10833_),
    .B2(_02574_),
    .C1(_10835_),
    .X(_03952_));
 sky130_fd_sc_hd__buf_1 _13592_ (.A(_10825_),
    .X(_10836_));
 sky130_fd_sc_hd__o221a_2 _13593_ (.A1(_10834_),
    .A2(\reg_pc[23] ),
    .B1(_10836_),
    .B2(_02573_),
    .C1(_10835_),
    .X(_03951_));
 sky130_fd_sc_hd__o221a_2 _13594_ (.A1(_10834_),
    .A2(\reg_pc[22] ),
    .B1(_10836_),
    .B2(_02572_),
    .C1(_10835_),
    .X(_03950_));
 sky130_fd_sc_hd__o221a_2 _13595_ (.A1(_10834_),
    .A2(\reg_pc[21] ),
    .B1(_10836_),
    .B2(_02570_),
    .C1(_10835_),
    .X(_03949_));
 sky130_fd_sc_hd__buf_1 _13596_ (.A(_10651_),
    .X(_10837_));
 sky130_fd_sc_hd__buf_1 _13597_ (.A(_10828_),
    .X(_10838_));
 sky130_fd_sc_hd__o221a_2 _13598_ (.A1(_10837_),
    .A2(\reg_pc[20] ),
    .B1(_10836_),
    .B2(_02569_),
    .C1(_10838_),
    .X(_03948_));
 sky130_fd_sc_hd__o221a_2 _13599_ (.A1(_10837_),
    .A2(\reg_pc[19] ),
    .B1(_10836_),
    .B2(_02568_),
    .C1(_10838_),
    .X(_03947_));
 sky130_fd_sc_hd__o221a_2 _13600_ (.A1(_10837_),
    .A2(\reg_pc[18] ),
    .B1(_10836_),
    .B2(_02567_),
    .C1(_10838_),
    .X(_03946_));
 sky130_fd_sc_hd__buf_1 _13601_ (.A(_10825_),
    .X(_10839_));
 sky130_fd_sc_hd__o221a_2 _13602_ (.A1(_10837_),
    .A2(\reg_pc[17] ),
    .B1(_10839_),
    .B2(_02566_),
    .C1(_10838_),
    .X(_03945_));
 sky130_fd_sc_hd__o221a_2 _13603_ (.A1(_10837_),
    .A2(\reg_pc[16] ),
    .B1(_10839_),
    .B2(_02565_),
    .C1(_10838_),
    .X(_03944_));
 sky130_fd_sc_hd__o221a_2 _13604_ (.A1(_10837_),
    .A2(\reg_pc[15] ),
    .B1(_10839_),
    .B2(_02564_),
    .C1(_10838_),
    .X(_03943_));
 sky130_fd_sc_hd__buf_1 _13605_ (.A(_10651_),
    .X(_10840_));
 sky130_fd_sc_hd__buf_1 _13606_ (.A(_10828_),
    .X(_10841_));
 sky130_fd_sc_hd__o221a_2 _13607_ (.A1(_10840_),
    .A2(\reg_pc[14] ),
    .B1(_10839_),
    .B2(_02563_),
    .C1(_10841_),
    .X(_03942_));
 sky130_fd_sc_hd__o221a_2 _13608_ (.A1(_10840_),
    .A2(\reg_pc[13] ),
    .B1(_10839_),
    .B2(_02562_),
    .C1(_10841_),
    .X(_03941_));
 sky130_fd_sc_hd__o221a_2 _13609_ (.A1(_10840_),
    .A2(\reg_pc[12] ),
    .B1(_10839_),
    .B2(_02561_),
    .C1(_10841_),
    .X(_03940_));
 sky130_fd_sc_hd__buf_1 _13610_ (.A(_10825_),
    .X(_10842_));
 sky130_fd_sc_hd__o221a_2 _13611_ (.A1(_10840_),
    .A2(\reg_pc[11] ),
    .B1(_10842_),
    .B2(_02589_),
    .C1(_10841_),
    .X(_03939_));
 sky130_fd_sc_hd__o221a_2 _13612_ (.A1(_10840_),
    .A2(\reg_pc[10] ),
    .B1(_10842_),
    .B2(_02588_),
    .C1(_10841_),
    .X(_03938_));
 sky130_fd_sc_hd__o221a_2 _13613_ (.A1(_10840_),
    .A2(\reg_pc[9] ),
    .B1(_10842_),
    .B2(_02587_),
    .C1(_10841_),
    .X(_03937_));
 sky130_fd_sc_hd__buf_1 _13614_ (.A(_10651_),
    .X(_10843_));
 sky130_fd_sc_hd__buf_1 _13615_ (.A(_10828_),
    .X(_10844_));
 sky130_fd_sc_hd__o221a_2 _13616_ (.A1(_10843_),
    .A2(\reg_pc[8] ),
    .B1(_10842_),
    .B2(_02586_),
    .C1(_10844_),
    .X(_03936_));
 sky130_fd_sc_hd__o221a_2 _13617_ (.A1(_10843_),
    .A2(\reg_pc[7] ),
    .B1(_10842_),
    .B2(_02585_),
    .C1(_10844_),
    .X(_03935_));
 sky130_fd_sc_hd__o221a_2 _13618_ (.A1(_10843_),
    .A2(\reg_pc[6] ),
    .B1(_10842_),
    .B2(_02584_),
    .C1(_10844_),
    .X(_03934_));
 sky130_fd_sc_hd__o221a_2 _13619_ (.A1(_10843_),
    .A2(\reg_pc[5] ),
    .B1(_10813_),
    .B2(_02583_),
    .C1(_10844_),
    .X(_03933_));
 sky130_fd_sc_hd__inv_2 _13620_ (.A(_01475_),
    .Y(_02582_));
 sky130_fd_sc_hd__o221a_2 _13621_ (.A1(_10843_),
    .A2(\reg_pc[4] ),
    .B1(_10813_),
    .B2(_02582_),
    .C1(_10844_),
    .X(_03932_));
 sky130_fd_sc_hd__o221a_2 _13622_ (.A1(_10843_),
    .A2(\reg_pc[3] ),
    .B1(_10813_),
    .B2(_02571_),
    .C1(_10844_),
    .X(_03931_));
 sky130_fd_sc_hd__buf_1 _13623_ (.A(_10444_),
    .X(_10845_));
 sky130_fd_sc_hd__buf_1 _13624_ (.A(_10845_),
    .X(_10846_));
 sky130_fd_sc_hd__o221a_2 _13625_ (.A1(_10652_),
    .A2(\reg_pc[2] ),
    .B1(_10813_),
    .B2(_02560_),
    .C1(_10846_),
    .X(_03930_));
 sky130_fd_sc_hd__o221a_2 _13626_ (.A1(_10652_),
    .A2(\reg_pc[1] ),
    .B1(_10813_),
    .B2(_02590_),
    .C1(_10846_),
    .X(_03929_));
 sky130_vsdinv _13627_ (.A(\count_instr[62] ),
    .Y(_10847_));
 sky130_vsdinv _13628_ (.A(\count_instr[61] ),
    .Y(_10848_));
 sky130_vsdinv _13629_ (.A(\count_instr[60] ),
    .Y(_10849_));
 sky130_vsdinv _13630_ (.A(\count_instr[59] ),
    .Y(_10850_));
 sky130_vsdinv _13631_ (.A(\count_instr[58] ),
    .Y(_10851_));
 sky130_vsdinv _13632_ (.A(\count_instr[57] ),
    .Y(_10852_));
 sky130_vsdinv _13633_ (.A(\count_instr[56] ),
    .Y(_10853_));
 sky130_vsdinv _13634_ (.A(\count_instr[55] ),
    .Y(_10854_));
 sky130_vsdinv _13635_ (.A(\count_instr[54] ),
    .Y(_10855_));
 sky130_vsdinv _13636_ (.A(\count_instr[53] ),
    .Y(_10856_));
 sky130_vsdinv _13637_ (.A(\count_instr[52] ),
    .Y(_10857_));
 sky130_vsdinv _13638_ (.A(\count_instr[51] ),
    .Y(_10858_));
 sky130_vsdinv _13639_ (.A(\count_instr[50] ),
    .Y(_10859_));
 sky130_vsdinv _13640_ (.A(\count_instr[49] ),
    .Y(_10860_));
 sky130_vsdinv _13641_ (.A(\count_instr[48] ),
    .Y(_10861_));
 sky130_vsdinv _13642_ (.A(\count_instr[47] ),
    .Y(_10862_));
 sky130_vsdinv _13643_ (.A(\count_instr[46] ),
    .Y(_10863_));
 sky130_vsdinv _13644_ (.A(\count_instr[45] ),
    .Y(_10864_));
 sky130_vsdinv _13645_ (.A(\count_instr[44] ),
    .Y(_10865_));
 sky130_vsdinv _13646_ (.A(\count_instr[43] ),
    .Y(_10866_));
 sky130_vsdinv _13647_ (.A(\count_instr[42] ),
    .Y(_10867_));
 sky130_vsdinv _13648_ (.A(\count_instr[41] ),
    .Y(_10868_));
 sky130_vsdinv _13649_ (.A(\count_instr[40] ),
    .Y(_10869_));
 sky130_vsdinv _13650_ (.A(\count_instr[39] ),
    .Y(_10870_));
 sky130_vsdinv _13651_ (.A(\count_instr[38] ),
    .Y(_10871_));
 sky130_vsdinv _13652_ (.A(\count_instr[37] ),
    .Y(_10872_));
 sky130_vsdinv _13653_ (.A(\count_instr[36] ),
    .Y(_10873_));
 sky130_vsdinv _13654_ (.A(\count_instr[35] ),
    .Y(_10874_));
 sky130_vsdinv _13655_ (.A(\count_instr[34] ),
    .Y(_10875_));
 sky130_vsdinv _13656_ (.A(\count_instr[33] ),
    .Y(_10876_));
 sky130_vsdinv _13657_ (.A(\count_instr[32] ),
    .Y(_10877_));
 sky130_vsdinv _13658_ (.A(\count_instr[31] ),
    .Y(_10878_));
 sky130_vsdinv _13659_ (.A(\count_instr[30] ),
    .Y(_10879_));
 sky130_vsdinv _13660_ (.A(\count_instr[29] ),
    .Y(_10880_));
 sky130_vsdinv _13661_ (.A(\count_instr[28] ),
    .Y(_10881_));
 sky130_vsdinv _13662_ (.A(\count_instr[27] ),
    .Y(_10882_));
 sky130_vsdinv _13663_ (.A(\count_instr[26] ),
    .Y(_10883_));
 sky130_vsdinv _13664_ (.A(\count_instr[25] ),
    .Y(_10884_));
 sky130_vsdinv _13665_ (.A(\count_instr[24] ),
    .Y(_10885_));
 sky130_vsdinv _13666_ (.A(\count_instr[23] ),
    .Y(_10886_));
 sky130_vsdinv _13667_ (.A(\count_instr[22] ),
    .Y(_10887_));
 sky130_vsdinv _13668_ (.A(\count_instr[21] ),
    .Y(_10888_));
 sky130_vsdinv _13669_ (.A(\count_instr[20] ),
    .Y(_10889_));
 sky130_vsdinv _13670_ (.A(\count_instr[19] ),
    .Y(_10890_));
 sky130_vsdinv _13671_ (.A(\count_instr[18] ),
    .Y(_10891_));
 sky130_vsdinv _13672_ (.A(\count_instr[17] ),
    .Y(_10892_));
 sky130_vsdinv _13673_ (.A(\count_instr[16] ),
    .Y(_10893_));
 sky130_vsdinv _13674_ (.A(\count_instr[15] ),
    .Y(_10894_));
 sky130_vsdinv _13675_ (.A(\count_instr[14] ),
    .Y(_10895_));
 sky130_vsdinv _13676_ (.A(\count_instr[13] ),
    .Y(_10896_));
 sky130_vsdinv _13677_ (.A(\count_instr[12] ),
    .Y(_10897_));
 sky130_vsdinv _13678_ (.A(\count_instr[11] ),
    .Y(_10898_));
 sky130_vsdinv _13679_ (.A(\count_instr[10] ),
    .Y(_10899_));
 sky130_vsdinv _13680_ (.A(\count_instr[9] ),
    .Y(_10900_));
 sky130_vsdinv _13681_ (.A(\count_instr[8] ),
    .Y(_10901_));
 sky130_vsdinv _13682_ (.A(\count_instr[7] ),
    .Y(_10902_));
 sky130_vsdinv _13683_ (.A(\count_instr[6] ),
    .Y(_10903_));
 sky130_vsdinv _13684_ (.A(\count_instr[5] ),
    .Y(_10904_));
 sky130_vsdinv _13685_ (.A(\count_instr[4] ),
    .Y(_10905_));
 sky130_vsdinv _13686_ (.A(\count_instr[3] ),
    .Y(_10906_));
 sky130_vsdinv _13687_ (.A(\count_instr[2] ),
    .Y(_10907_));
 sky130_vsdinv _13688_ (.A(\count_instr[1] ),
    .Y(_10908_));
 sky130_vsdinv _13689_ (.A(\count_instr[0] ),
    .Y(_10909_));
 sky130_fd_sc_hd__or2_2 _13690_ (.A(_10909_),
    .B(_10566_),
    .X(_10910_));
 sky130_fd_sc_hd__or3_2 _13691_ (.A(_10907_),
    .B(_10908_),
    .C(_10910_),
    .X(_10911_));
 sky130_fd_sc_hd__or2_2 _13692_ (.A(_10906_),
    .B(_10911_),
    .X(_10912_));
 sky130_fd_sc_hd__or2_2 _13693_ (.A(_10905_),
    .B(_10912_),
    .X(_10913_));
 sky130_fd_sc_hd__or2_2 _13694_ (.A(_10904_),
    .B(_10913_),
    .X(_10914_));
 sky130_fd_sc_hd__or2_2 _13695_ (.A(_10903_),
    .B(_10914_),
    .X(_10915_));
 sky130_fd_sc_hd__or2_2 _13696_ (.A(_10902_),
    .B(_10915_),
    .X(_10916_));
 sky130_fd_sc_hd__or2_2 _13697_ (.A(_10901_),
    .B(_10916_),
    .X(_10917_));
 sky130_fd_sc_hd__or2_2 _13698_ (.A(_10900_),
    .B(_10917_),
    .X(_10918_));
 sky130_fd_sc_hd__or2_2 _13699_ (.A(_10899_),
    .B(_10918_),
    .X(_10919_));
 sky130_fd_sc_hd__or2_2 _13700_ (.A(_10898_),
    .B(_10919_),
    .X(_10920_));
 sky130_fd_sc_hd__or2_2 _13701_ (.A(_10897_),
    .B(_10920_),
    .X(_10921_));
 sky130_fd_sc_hd__or2_2 _13702_ (.A(_10896_),
    .B(_10921_),
    .X(_10922_));
 sky130_fd_sc_hd__or2_2 _13703_ (.A(_10895_),
    .B(_10922_),
    .X(_10923_));
 sky130_fd_sc_hd__or2_2 _13704_ (.A(_10894_),
    .B(_10923_),
    .X(_10924_));
 sky130_fd_sc_hd__or2_2 _13705_ (.A(_10893_),
    .B(_10924_),
    .X(_10925_));
 sky130_fd_sc_hd__or2_2 _13706_ (.A(_10892_),
    .B(_10925_),
    .X(_10926_));
 sky130_fd_sc_hd__or2_2 _13707_ (.A(_10891_),
    .B(_10926_),
    .X(_10927_));
 sky130_fd_sc_hd__or2_2 _13708_ (.A(_10890_),
    .B(_10927_),
    .X(_10928_));
 sky130_fd_sc_hd__or2_2 _13709_ (.A(_10889_),
    .B(_10928_),
    .X(_10929_));
 sky130_fd_sc_hd__or2_2 _13710_ (.A(_10888_),
    .B(_10929_),
    .X(_10930_));
 sky130_fd_sc_hd__or2_2 _13711_ (.A(_10887_),
    .B(_10930_),
    .X(_10931_));
 sky130_fd_sc_hd__or2_2 _13712_ (.A(_10886_),
    .B(_10931_),
    .X(_10932_));
 sky130_fd_sc_hd__or2_2 _13713_ (.A(_10885_),
    .B(_10932_),
    .X(_10933_));
 sky130_fd_sc_hd__or2_2 _13714_ (.A(_10884_),
    .B(_10933_),
    .X(_10934_));
 sky130_fd_sc_hd__or2_2 _13715_ (.A(_10883_),
    .B(_10934_),
    .X(_10935_));
 sky130_fd_sc_hd__or2_2 _13716_ (.A(_10882_),
    .B(_10935_),
    .X(_10936_));
 sky130_fd_sc_hd__or2_2 _13717_ (.A(_10881_),
    .B(_10936_),
    .X(_10937_));
 sky130_fd_sc_hd__or2_2 _13718_ (.A(_10880_),
    .B(_10937_),
    .X(_10938_));
 sky130_fd_sc_hd__or2_2 _13719_ (.A(_10879_),
    .B(_10938_),
    .X(_10939_));
 sky130_fd_sc_hd__or2_2 _13720_ (.A(_10878_),
    .B(_10939_),
    .X(_10940_));
 sky130_fd_sc_hd__or2_2 _13721_ (.A(_10877_),
    .B(_10940_),
    .X(_10941_));
 sky130_fd_sc_hd__or2_2 _13722_ (.A(_10876_),
    .B(_10941_),
    .X(_10942_));
 sky130_fd_sc_hd__or2_2 _13723_ (.A(_10875_),
    .B(_10942_),
    .X(_10943_));
 sky130_fd_sc_hd__or2_2 _13724_ (.A(_10874_),
    .B(_10943_),
    .X(_10944_));
 sky130_fd_sc_hd__or2_2 _13725_ (.A(_10873_),
    .B(_10944_),
    .X(_10945_));
 sky130_fd_sc_hd__or2_2 _13726_ (.A(_10872_),
    .B(_10945_),
    .X(_10946_));
 sky130_fd_sc_hd__or2_2 _13727_ (.A(_10871_),
    .B(_10946_),
    .X(_10947_));
 sky130_fd_sc_hd__or2_2 _13728_ (.A(_10870_),
    .B(_10947_),
    .X(_10948_));
 sky130_fd_sc_hd__or2_2 _13729_ (.A(_10869_),
    .B(_10948_),
    .X(_10949_));
 sky130_fd_sc_hd__or2_2 _13730_ (.A(_10868_),
    .B(_10949_),
    .X(_10950_));
 sky130_fd_sc_hd__or2_2 _13731_ (.A(_10867_),
    .B(_10950_),
    .X(_10951_));
 sky130_fd_sc_hd__or2_2 _13732_ (.A(_10866_),
    .B(_10951_),
    .X(_10952_));
 sky130_fd_sc_hd__or2_2 _13733_ (.A(_10865_),
    .B(_10952_),
    .X(_10953_));
 sky130_fd_sc_hd__or2_2 _13734_ (.A(_10864_),
    .B(_10953_),
    .X(_10954_));
 sky130_fd_sc_hd__or2_2 _13735_ (.A(_10863_),
    .B(_10954_),
    .X(_10955_));
 sky130_fd_sc_hd__or2_2 _13736_ (.A(_10862_),
    .B(_10955_),
    .X(_10956_));
 sky130_fd_sc_hd__or2_2 _13737_ (.A(_10861_),
    .B(_10956_),
    .X(_10957_));
 sky130_fd_sc_hd__or2_2 _13738_ (.A(_10860_),
    .B(_10957_),
    .X(_10958_));
 sky130_fd_sc_hd__or2_2 _13739_ (.A(_10859_),
    .B(_10958_),
    .X(_10959_));
 sky130_fd_sc_hd__or2_2 _13740_ (.A(_10858_),
    .B(_10959_),
    .X(_10960_));
 sky130_fd_sc_hd__or2_2 _13741_ (.A(_10857_),
    .B(_10960_),
    .X(_10961_));
 sky130_fd_sc_hd__or2_2 _13742_ (.A(_10856_),
    .B(_10961_),
    .X(_10962_));
 sky130_fd_sc_hd__or2_2 _13743_ (.A(_10855_),
    .B(_10962_),
    .X(_10963_));
 sky130_fd_sc_hd__or2_2 _13744_ (.A(_10854_),
    .B(_10963_),
    .X(_10964_));
 sky130_fd_sc_hd__or2_2 _13745_ (.A(_10853_),
    .B(_10964_),
    .X(_10965_));
 sky130_fd_sc_hd__or2_2 _13746_ (.A(_10852_),
    .B(_10965_),
    .X(_10966_));
 sky130_fd_sc_hd__or2_2 _13747_ (.A(_10851_),
    .B(_10966_),
    .X(_10967_));
 sky130_fd_sc_hd__or2_2 _13748_ (.A(_10850_),
    .B(_10967_),
    .X(_10968_));
 sky130_fd_sc_hd__or2_2 _13749_ (.A(_10849_),
    .B(_10968_),
    .X(_10969_));
 sky130_fd_sc_hd__or2_2 _13750_ (.A(_10848_),
    .B(_10969_),
    .X(_10970_));
 sky130_fd_sc_hd__or2_2 _13751_ (.A(_10847_),
    .B(_10970_),
    .X(_10971_));
 sky130_vsdinv _13752_ (.A(_10971_),
    .Y(_10972_));
 sky130_vsdinv _13753_ (.A(\count_instr[63] ),
    .Y(_10973_));
 sky130_fd_sc_hd__o221a_2 _13754_ (.A1(\count_instr[63] ),
    .A2(_10972_),
    .B1(_10973_),
    .B2(_10971_),
    .C1(_10846_),
    .X(_03928_));
 sky130_fd_sc_hd__buf_1 _13755_ (.A(_10688_),
    .X(_10974_));
 sky130_fd_sc_hd__a211oi_2 _13756_ (.A1(_10847_),
    .A2(_10970_),
    .B1(_10974_),
    .C1(_10972_),
    .Y(_03927_));
 sky130_vsdinv _13757_ (.A(_10969_),
    .Y(_10975_));
 sky130_fd_sc_hd__o211a_2 _13758_ (.A1(\count_instr[61] ),
    .A2(_10975_),
    .B1(_10658_),
    .C1(_10970_),
    .X(_03926_));
 sky130_fd_sc_hd__a211oi_2 _13759_ (.A1(_10849_),
    .A2(_10968_),
    .B1(_10974_),
    .C1(_10975_),
    .Y(_03925_));
 sky130_vsdinv _13760_ (.A(_10967_),
    .Y(_10976_));
 sky130_fd_sc_hd__o211a_2 _13761_ (.A1(\count_instr[59] ),
    .A2(_10976_),
    .B1(_10658_),
    .C1(_10968_),
    .X(_03924_));
 sky130_fd_sc_hd__a211oi_2 _13762_ (.A1(_10851_),
    .A2(_10966_),
    .B1(_10974_),
    .C1(_10976_),
    .Y(_03923_));
 sky130_vsdinv _13763_ (.A(_10965_),
    .Y(_10977_));
 sky130_fd_sc_hd__o211a_2 _13764_ (.A1(\count_instr[57] ),
    .A2(_10977_),
    .B1(_10658_),
    .C1(_10966_),
    .X(_03922_));
 sky130_fd_sc_hd__a211oi_2 _13765_ (.A1(_10853_),
    .A2(_10964_),
    .B1(_10974_),
    .C1(_10977_),
    .Y(_03921_));
 sky130_vsdinv _13766_ (.A(_10963_),
    .Y(_10978_));
 sky130_fd_sc_hd__o211a_2 _13767_ (.A1(\count_instr[55] ),
    .A2(_10978_),
    .B1(_10658_),
    .C1(_10964_),
    .X(_03920_));
 sky130_fd_sc_hd__a211oi_2 _13768_ (.A1(_10855_),
    .A2(_10962_),
    .B1(_10974_),
    .C1(_10978_),
    .Y(_03919_));
 sky130_vsdinv _13769_ (.A(_10961_),
    .Y(_10979_));
 sky130_fd_sc_hd__o211a_2 _13770_ (.A1(\count_instr[53] ),
    .A2(_10979_),
    .B1(_10658_),
    .C1(_10962_),
    .X(_03918_));
 sky130_fd_sc_hd__buf_1 _13771_ (.A(_10774_),
    .X(_10980_));
 sky130_fd_sc_hd__a211oi_2 _13772_ (.A1(_10857_),
    .A2(_10960_),
    .B1(_10980_),
    .C1(_10979_),
    .Y(_03917_));
 sky130_vsdinv _13773_ (.A(_10959_),
    .Y(_10981_));
 sky130_fd_sc_hd__buf_1 _13774_ (.A(_10463_),
    .X(_10982_));
 sky130_fd_sc_hd__o211a_2 _13775_ (.A1(\count_instr[51] ),
    .A2(_10981_),
    .B1(_10982_),
    .C1(_10960_),
    .X(_03916_));
 sky130_fd_sc_hd__a211oi_2 _13776_ (.A1(_10859_),
    .A2(_10958_),
    .B1(_10980_),
    .C1(_10981_),
    .Y(_03915_));
 sky130_vsdinv _13777_ (.A(_10957_),
    .Y(_10983_));
 sky130_fd_sc_hd__o211a_2 _13778_ (.A1(\count_instr[49] ),
    .A2(_10983_),
    .B1(_10982_),
    .C1(_10958_),
    .X(_03914_));
 sky130_fd_sc_hd__a211oi_2 _13779_ (.A1(_10861_),
    .A2(_10956_),
    .B1(_10980_),
    .C1(_10983_),
    .Y(_03913_));
 sky130_vsdinv _13780_ (.A(_10955_),
    .Y(_10984_));
 sky130_fd_sc_hd__o211a_2 _13781_ (.A1(\count_instr[47] ),
    .A2(_10984_),
    .B1(_10982_),
    .C1(_10956_),
    .X(_03912_));
 sky130_fd_sc_hd__a211oi_2 _13782_ (.A1(_10863_),
    .A2(_10954_),
    .B1(_10980_),
    .C1(_10984_),
    .Y(_03911_));
 sky130_vsdinv _13783_ (.A(_10953_),
    .Y(_10985_));
 sky130_fd_sc_hd__o211a_2 _13784_ (.A1(\count_instr[45] ),
    .A2(_10985_),
    .B1(_10982_),
    .C1(_10954_),
    .X(_03910_));
 sky130_fd_sc_hd__a211oi_2 _13785_ (.A1(_10865_),
    .A2(_10952_),
    .B1(_10980_),
    .C1(_10985_),
    .Y(_03909_));
 sky130_vsdinv _13786_ (.A(_10951_),
    .Y(_10986_));
 sky130_fd_sc_hd__o211a_2 _13787_ (.A1(\count_instr[43] ),
    .A2(_10986_),
    .B1(_10982_),
    .C1(_10952_),
    .X(_03908_));
 sky130_fd_sc_hd__a211oi_2 _13788_ (.A1(_10867_),
    .A2(_10950_),
    .B1(_10980_),
    .C1(_10986_),
    .Y(_03907_));
 sky130_vsdinv _13789_ (.A(_10949_),
    .Y(_10987_));
 sky130_fd_sc_hd__o211a_2 _13790_ (.A1(\count_instr[41] ),
    .A2(_10987_),
    .B1(_10982_),
    .C1(_10950_),
    .X(_03906_));
 sky130_fd_sc_hd__buf_1 _13791_ (.A(_10774_),
    .X(_10988_));
 sky130_fd_sc_hd__a211oi_2 _13792_ (.A1(_10869_),
    .A2(_10948_),
    .B1(_10988_),
    .C1(_10987_),
    .Y(_03905_));
 sky130_vsdinv _13793_ (.A(_10947_),
    .Y(_10989_));
 sky130_fd_sc_hd__buf_1 _13794_ (.A(_10463_),
    .X(_10990_));
 sky130_fd_sc_hd__o211a_2 _13795_ (.A1(\count_instr[39] ),
    .A2(_10989_),
    .B1(_10990_),
    .C1(_10948_),
    .X(_03904_));
 sky130_fd_sc_hd__a211oi_2 _13796_ (.A1(_10871_),
    .A2(_10946_),
    .B1(_10988_),
    .C1(_10989_),
    .Y(_03903_));
 sky130_vsdinv _13797_ (.A(_10945_),
    .Y(_10991_));
 sky130_fd_sc_hd__o211a_2 _13798_ (.A1(\count_instr[37] ),
    .A2(_10991_),
    .B1(_10990_),
    .C1(_10946_),
    .X(_03902_));
 sky130_fd_sc_hd__a211oi_2 _13799_ (.A1(_10873_),
    .A2(_10944_),
    .B1(_10988_),
    .C1(_10991_),
    .Y(_03901_));
 sky130_vsdinv _13800_ (.A(_10943_),
    .Y(_10992_));
 sky130_fd_sc_hd__o211a_2 _13801_ (.A1(\count_instr[35] ),
    .A2(_10992_),
    .B1(_10990_),
    .C1(_10944_),
    .X(_03900_));
 sky130_fd_sc_hd__a211oi_2 _13802_ (.A1(_10875_),
    .A2(_10942_),
    .B1(_10988_),
    .C1(_10992_),
    .Y(_03899_));
 sky130_vsdinv _13803_ (.A(_10941_),
    .Y(_10993_));
 sky130_fd_sc_hd__o211a_2 _13804_ (.A1(\count_instr[33] ),
    .A2(_10993_),
    .B1(_10990_),
    .C1(_10942_),
    .X(_03898_));
 sky130_fd_sc_hd__a211oi_2 _13805_ (.A1(_10877_),
    .A2(_10940_),
    .B1(_10988_),
    .C1(_10993_),
    .Y(_03897_));
 sky130_vsdinv _13806_ (.A(_10939_),
    .Y(_10994_));
 sky130_fd_sc_hd__o211a_2 _13807_ (.A1(\count_instr[31] ),
    .A2(_10994_),
    .B1(_10990_),
    .C1(_10940_),
    .X(_03896_));
 sky130_fd_sc_hd__a211oi_2 _13808_ (.A1(_10879_),
    .A2(_10938_),
    .B1(_10988_),
    .C1(_10994_),
    .Y(_03895_));
 sky130_vsdinv _13809_ (.A(_10937_),
    .Y(_10995_));
 sky130_fd_sc_hd__o211a_2 _13810_ (.A1(\count_instr[29] ),
    .A2(_10995_),
    .B1(_10990_),
    .C1(_10938_),
    .X(_03894_));
 sky130_fd_sc_hd__buf_1 _13811_ (.A(_10481_),
    .X(_10996_));
 sky130_fd_sc_hd__buf_1 _13812_ (.A(_10996_),
    .X(_10997_));
 sky130_fd_sc_hd__a211oi_2 _13813_ (.A1(_10881_),
    .A2(_10936_),
    .B1(_10997_),
    .C1(_10995_),
    .Y(_03893_));
 sky130_vsdinv _13814_ (.A(_10935_),
    .Y(_10998_));
 sky130_fd_sc_hd__buf_1 _13815_ (.A(_10463_),
    .X(_10999_));
 sky130_fd_sc_hd__o211a_2 _13816_ (.A1(\count_instr[27] ),
    .A2(_10998_),
    .B1(_10999_),
    .C1(_10936_),
    .X(_03892_));
 sky130_fd_sc_hd__a211oi_2 _13817_ (.A1(_10883_),
    .A2(_10934_),
    .B1(_10997_),
    .C1(_10998_),
    .Y(_03891_));
 sky130_vsdinv _13818_ (.A(_10933_),
    .Y(_11000_));
 sky130_fd_sc_hd__o211a_2 _13819_ (.A1(\count_instr[25] ),
    .A2(_11000_),
    .B1(_10999_),
    .C1(_10934_),
    .X(_03890_));
 sky130_fd_sc_hd__a211oi_2 _13820_ (.A1(_10885_),
    .A2(_10932_),
    .B1(_10997_),
    .C1(_11000_),
    .Y(_03889_));
 sky130_vsdinv _13821_ (.A(_10931_),
    .Y(_11001_));
 sky130_fd_sc_hd__o211a_2 _13822_ (.A1(\count_instr[23] ),
    .A2(_11001_),
    .B1(_10999_),
    .C1(_10932_),
    .X(_03888_));
 sky130_fd_sc_hd__a211oi_2 _13823_ (.A1(_10887_),
    .A2(_10930_),
    .B1(_10997_),
    .C1(_11001_),
    .Y(_03887_));
 sky130_vsdinv _13824_ (.A(_10929_),
    .Y(_11002_));
 sky130_fd_sc_hd__o211a_2 _13825_ (.A1(\count_instr[21] ),
    .A2(_11002_),
    .B1(_10999_),
    .C1(_10930_),
    .X(_03886_));
 sky130_fd_sc_hd__a211oi_2 _13826_ (.A1(_10889_),
    .A2(_10928_),
    .B1(_10997_),
    .C1(_11002_),
    .Y(_03885_));
 sky130_vsdinv _13827_ (.A(_10927_),
    .Y(_11003_));
 sky130_fd_sc_hd__o211a_2 _13828_ (.A1(\count_instr[19] ),
    .A2(_11003_),
    .B1(_10999_),
    .C1(_10928_),
    .X(_03884_));
 sky130_fd_sc_hd__a211oi_2 _13829_ (.A1(_10891_),
    .A2(_10926_),
    .B1(_10997_),
    .C1(_11003_),
    .Y(_03883_));
 sky130_vsdinv _13830_ (.A(_10925_),
    .Y(_11004_));
 sky130_fd_sc_hd__o211a_2 _13831_ (.A1(\count_instr[17] ),
    .A2(_11004_),
    .B1(_10999_),
    .C1(_10926_),
    .X(_03882_));
 sky130_fd_sc_hd__buf_1 _13832_ (.A(_10996_),
    .X(_11005_));
 sky130_fd_sc_hd__a211oi_2 _13833_ (.A1(_10893_),
    .A2(_10924_),
    .B1(_11005_),
    .C1(_11004_),
    .Y(_03881_));
 sky130_vsdinv _13834_ (.A(_10923_),
    .Y(_11006_));
 sky130_fd_sc_hd__buf_1 _13835_ (.A(_10443_),
    .X(_11007_));
 sky130_fd_sc_hd__buf_1 _13836_ (.A(_11007_),
    .X(_11008_));
 sky130_fd_sc_hd__o211a_2 _13837_ (.A1(\count_instr[15] ),
    .A2(_11006_),
    .B1(_11008_),
    .C1(_10924_),
    .X(_03880_));
 sky130_fd_sc_hd__a211oi_2 _13838_ (.A1(_10895_),
    .A2(_10922_),
    .B1(_11005_),
    .C1(_11006_),
    .Y(_03879_));
 sky130_vsdinv _13839_ (.A(_10921_),
    .Y(_11009_));
 sky130_fd_sc_hd__o211a_2 _13840_ (.A1(\count_instr[13] ),
    .A2(_11009_),
    .B1(_11008_),
    .C1(_10922_),
    .X(_03878_));
 sky130_fd_sc_hd__a211oi_2 _13841_ (.A1(_10897_),
    .A2(_10920_),
    .B1(_11005_),
    .C1(_11009_),
    .Y(_03877_));
 sky130_vsdinv _13842_ (.A(_10919_),
    .Y(_11010_));
 sky130_fd_sc_hd__o211a_2 _13843_ (.A1(\count_instr[11] ),
    .A2(_11010_),
    .B1(_11008_),
    .C1(_10920_),
    .X(_03876_));
 sky130_fd_sc_hd__a211oi_2 _13844_ (.A1(_10899_),
    .A2(_10918_),
    .B1(_11005_),
    .C1(_11010_),
    .Y(_03875_));
 sky130_vsdinv _13845_ (.A(_10917_),
    .Y(_11011_));
 sky130_fd_sc_hd__o211a_2 _13846_ (.A1(\count_instr[9] ),
    .A2(_11011_),
    .B1(_11008_),
    .C1(_10918_),
    .X(_03874_));
 sky130_fd_sc_hd__a211oi_2 _13847_ (.A1(_10901_),
    .A2(_10916_),
    .B1(_11005_),
    .C1(_11011_),
    .Y(_03873_));
 sky130_vsdinv _13848_ (.A(_10915_),
    .Y(_11012_));
 sky130_fd_sc_hd__o211a_2 _13849_ (.A1(\count_instr[7] ),
    .A2(_11012_),
    .B1(_11008_),
    .C1(_10916_),
    .X(_03872_));
 sky130_fd_sc_hd__a211oi_2 _13850_ (.A1(_10903_),
    .A2(_10914_),
    .B1(_11005_),
    .C1(_11012_),
    .Y(_03871_));
 sky130_vsdinv _13851_ (.A(_10913_),
    .Y(_11013_));
 sky130_fd_sc_hd__o211a_2 _13852_ (.A1(\count_instr[5] ),
    .A2(_11013_),
    .B1(_11008_),
    .C1(_10914_),
    .X(_03870_));
 sky130_fd_sc_hd__buf_1 _13853_ (.A(_10996_),
    .X(_11014_));
 sky130_fd_sc_hd__a211oi_2 _13854_ (.A1(_10905_),
    .A2(_10912_),
    .B1(_11014_),
    .C1(_11013_),
    .Y(_03869_));
 sky130_vsdinv _13855_ (.A(_10911_),
    .Y(_11015_));
 sky130_fd_sc_hd__buf_1 _13856_ (.A(_11007_),
    .X(_11016_));
 sky130_fd_sc_hd__o211a_2 _13857_ (.A1(\count_instr[3] ),
    .A2(_11015_),
    .B1(_11016_),
    .C1(_10912_),
    .X(_03868_));
 sky130_fd_sc_hd__buf_1 _13858_ (.A(_10774_),
    .X(_11017_));
 sky130_fd_sc_hd__o21a_2 _13859_ (.A1(_10908_),
    .A2(_10910_),
    .B1(_10907_),
    .X(_11018_));
 sky130_fd_sc_hd__nor3_2 _13860_ (.A(_11017_),
    .B(_11015_),
    .C(_11018_),
    .Y(_03867_));
 sky130_vsdinv _13861_ (.A(_10910_),
    .Y(_11019_));
 sky130_fd_sc_hd__o221a_2 _13862_ (.A1(_10908_),
    .A2(_10910_),
    .B1(\count_instr[1] ),
    .B2(_11019_),
    .C1(_10846_),
    .X(_03866_));
 sky130_fd_sc_hd__o211a_2 _13863_ (.A1(\count_instr[0] ),
    .A2(_10567_),
    .B1(_11016_),
    .C1(_10910_),
    .X(_03865_));
 sky130_fd_sc_hd__or2_2 _13864_ (.A(\cpu_state[1] ),
    .B(\cpu_state[2] ),
    .X(_11020_));
 sky130_fd_sc_hd__o221a_2 _13865_ (.A1(instr_retirq),
    .A2(_10468_),
    .B1(\irq_state[1] ),
    .B2(_10508_),
    .C1(_11020_),
    .X(_11021_));
 sky130_fd_sc_hd__buf_1 _13866_ (.A(_11021_),
    .X(_11022_));
 sky130_fd_sc_hd__buf_1 _13867_ (.A(_11022_),
    .X(_11023_));
 sky130_vsdinv _13868_ (.A(_11021_),
    .Y(_11024_));
 sky130_fd_sc_hd__buf_1 _13869_ (.A(_11024_),
    .X(_11025_));
 sky130_fd_sc_hd__buf_1 _13870_ (.A(_11025_),
    .X(_11026_));
 sky130_fd_sc_hd__buf_1 _13871_ (.A(_10614_),
    .X(_11027_));
 sky130_fd_sc_hd__buf_1 _13872_ (.A(_11027_),
    .X(_11028_));
 sky130_fd_sc_hd__nor3_2 _13873_ (.A(\irq_mask[31] ),
    .B(_10544_),
    .C(_11028_),
    .Y(_11029_));
 sky130_fd_sc_hd__o221a_2 _13874_ (.A1(eoi[31]),
    .A2(_11023_),
    .B1(_11026_),
    .B2(_11029_),
    .C1(_10846_),
    .X(_03864_));
 sky130_fd_sc_hd__buf_1 _13875_ (.A(_10469_),
    .X(_11030_));
 sky130_fd_sc_hd__buf_1 _13876_ (.A(_11030_),
    .X(_11031_));
 sky130_fd_sc_hd__and3_2 _13877_ (.A(_10542_),
    .B(\irq_pending[30] ),
    .C(_11031_),
    .X(_11032_));
 sky130_fd_sc_hd__o221a_2 _13878_ (.A1(eoi[30]),
    .A2(_11023_),
    .B1(_11026_),
    .B2(_11032_),
    .C1(_10846_),
    .X(_03863_));
 sky130_fd_sc_hd__nor3_2 _13879_ (.A(\irq_mask[29] ),
    .B(_10543_),
    .C(_11028_),
    .Y(_11033_));
 sky130_fd_sc_hd__buf_1 _13880_ (.A(_10845_),
    .X(_11034_));
 sky130_fd_sc_hd__o221a_2 _13881_ (.A1(eoi[29]),
    .A2(_11023_),
    .B1(_11026_),
    .B2(_11033_),
    .C1(_11034_),
    .X(_03862_));
 sky130_fd_sc_hd__and3_2 _13882_ (.A(_10541_),
    .B(\irq_pending[28] ),
    .C(_11031_),
    .X(_11035_));
 sky130_fd_sc_hd__o221a_2 _13883_ (.A1(eoi[28]),
    .A2(_11023_),
    .B1(_11026_),
    .B2(_11035_),
    .C1(_11034_),
    .X(_03861_));
 sky130_fd_sc_hd__nor3_2 _13884_ (.A(\irq_mask[27] ),
    .B(_10525_),
    .C(_11028_),
    .Y(_11036_));
 sky130_fd_sc_hd__o221a_2 _13885_ (.A1(eoi[27]),
    .A2(_11023_),
    .B1(_11026_),
    .B2(_11036_),
    .C1(_11034_),
    .X(_03860_));
 sky130_fd_sc_hd__and3_2 _13886_ (.A(_10523_),
    .B(\irq_pending[26] ),
    .C(_11031_),
    .X(_11037_));
 sky130_fd_sc_hd__o221a_2 _13887_ (.A1(eoi[26]),
    .A2(_11023_),
    .B1(_11026_),
    .B2(_11037_),
    .C1(_11034_),
    .X(_03859_));
 sky130_fd_sc_hd__buf_1 _13888_ (.A(_11022_),
    .X(_11038_));
 sky130_fd_sc_hd__buf_1 _13889_ (.A(_11025_),
    .X(_11039_));
 sky130_fd_sc_hd__nor3_2 _13890_ (.A(\irq_mask[25] ),
    .B(_10524_),
    .C(_11028_),
    .Y(_11040_));
 sky130_fd_sc_hd__o221a_2 _13891_ (.A1(eoi[25]),
    .A2(_11038_),
    .B1(_11039_),
    .B2(_11040_),
    .C1(_11034_),
    .X(_03858_));
 sky130_fd_sc_hd__buf_1 _13892_ (.A(_11030_),
    .X(_11041_));
 sky130_fd_sc_hd__and3_2 _13893_ (.A(_10522_),
    .B(\irq_pending[24] ),
    .C(_11041_),
    .X(_11042_));
 sky130_fd_sc_hd__o221a_2 _13894_ (.A1(eoi[24]),
    .A2(_11038_),
    .B1(_11039_),
    .B2(_11042_),
    .C1(_11034_),
    .X(_03857_));
 sky130_fd_sc_hd__nor3_2 _13895_ (.A(\irq_mask[23] ),
    .B(_10556_),
    .C(_11028_),
    .Y(_11043_));
 sky130_fd_sc_hd__buf_1 _13896_ (.A(_10845_),
    .X(_11044_));
 sky130_fd_sc_hd__o221a_2 _13897_ (.A1(eoi[23]),
    .A2(_11038_),
    .B1(_11039_),
    .B2(_11043_),
    .C1(_11044_),
    .X(_03856_));
 sky130_fd_sc_hd__and3_2 _13898_ (.A(_10554_),
    .B(\irq_pending[22] ),
    .C(_11041_),
    .X(_11045_));
 sky130_fd_sc_hd__o221a_2 _13899_ (.A1(eoi[22]),
    .A2(_11038_),
    .B1(_11039_),
    .B2(_11045_),
    .C1(_11044_),
    .X(_03855_));
 sky130_fd_sc_hd__nor3_2 _13900_ (.A(\irq_mask[21] ),
    .B(_10555_),
    .C(_11028_),
    .Y(_11046_));
 sky130_fd_sc_hd__o221a_2 _13901_ (.A1(eoi[21]),
    .A2(_11038_),
    .B1(_11039_),
    .B2(_11046_),
    .C1(_11044_),
    .X(_03854_));
 sky130_fd_sc_hd__and3_2 _13902_ (.A(_10553_),
    .B(\irq_pending[20] ),
    .C(_11041_),
    .X(_11047_));
 sky130_fd_sc_hd__o221a_2 _13903_ (.A1(eoi[20]),
    .A2(_11038_),
    .B1(_11039_),
    .B2(_11047_),
    .C1(_11044_),
    .X(_03853_));
 sky130_fd_sc_hd__buf_1 _13904_ (.A(_11022_),
    .X(_11048_));
 sky130_fd_sc_hd__buf_1 _13905_ (.A(_11025_),
    .X(_11049_));
 sky130_fd_sc_hd__buf_1 _13906_ (.A(_10614_),
    .X(_11050_));
 sky130_fd_sc_hd__nor3_2 _13907_ (.A(\irq_mask[19] ),
    .B(_10517_),
    .C(_11050_),
    .Y(_11051_));
 sky130_fd_sc_hd__o221a_2 _13908_ (.A1(eoi[19]),
    .A2(_11048_),
    .B1(_11049_),
    .B2(_11051_),
    .C1(_11044_),
    .X(_03852_));
 sky130_vsdinv _13909_ (.A(\irq_mask[18] ),
    .Y(_11052_));
 sky130_fd_sc_hd__and3_2 _13910_ (.A(_11052_),
    .B(\irq_pending[18] ),
    .C(_11041_),
    .X(_11053_));
 sky130_fd_sc_hd__o221a_2 _13911_ (.A1(eoi[18]),
    .A2(_11048_),
    .B1(_11049_),
    .B2(_11053_),
    .C1(_11044_),
    .X(_03851_));
 sky130_fd_sc_hd__nor3_2 _13912_ (.A(\irq_mask[17] ),
    .B(_10516_),
    .C(_11050_),
    .Y(_11054_));
 sky130_fd_sc_hd__buf_1 _13913_ (.A(_10845_),
    .X(_11055_));
 sky130_fd_sc_hd__o221a_2 _13914_ (.A1(eoi[17]),
    .A2(_11048_),
    .B1(_11049_),
    .B2(_11054_),
    .C1(_11055_),
    .X(_03850_));
 sky130_fd_sc_hd__nor3_2 _13915_ (.A(\irq_mask[16] ),
    .B(_10518_),
    .C(_11050_),
    .Y(_11056_));
 sky130_fd_sc_hd__o221a_2 _13916_ (.A1(eoi[16]),
    .A2(_11048_),
    .B1(_11049_),
    .B2(_11056_),
    .C1(_11055_),
    .X(_03849_));
 sky130_fd_sc_hd__and3_2 _13917_ (.A(_10536_),
    .B(\irq_pending[15] ),
    .C(_11041_),
    .X(_11057_));
 sky130_fd_sc_hd__o221a_2 _13918_ (.A1(eoi[15]),
    .A2(_11048_),
    .B1(_11049_),
    .B2(_11057_),
    .C1(_11055_),
    .X(_03848_));
 sky130_fd_sc_hd__nor3_2 _13919_ (.A(\irq_mask[14] ),
    .B(_10538_),
    .C(_11050_),
    .Y(_11058_));
 sky130_fd_sc_hd__o221a_2 _13920_ (.A1(eoi[14]),
    .A2(_11048_),
    .B1(_11049_),
    .B2(_11058_),
    .C1(_11055_),
    .X(_03847_));
 sky130_fd_sc_hd__buf_1 _13921_ (.A(_11022_),
    .X(_11059_));
 sky130_fd_sc_hd__buf_1 _13922_ (.A(_11025_),
    .X(_11060_));
 sky130_fd_sc_hd__and3_2 _13923_ (.A(_10535_),
    .B(\irq_pending[13] ),
    .C(_11041_),
    .X(_11061_));
 sky130_fd_sc_hd__o221a_2 _13924_ (.A1(eoi[13]),
    .A2(_11059_),
    .B1(_11060_),
    .B2(_11061_),
    .C1(_11055_),
    .X(_03846_));
 sky130_fd_sc_hd__nor3_2 _13925_ (.A(\irq_mask[12] ),
    .B(_10537_),
    .C(_11050_),
    .Y(_11062_));
 sky130_fd_sc_hd__o221a_2 _13926_ (.A1(eoi[12]),
    .A2(_11059_),
    .B1(_11060_),
    .B2(_11062_),
    .C1(_11055_),
    .X(_03845_));
 sky130_fd_sc_hd__buf_1 _13927_ (.A(_11030_),
    .X(_11063_));
 sky130_fd_sc_hd__and3_2 _13928_ (.A(_10548_),
    .B(\irq_pending[11] ),
    .C(_11063_),
    .X(_11064_));
 sky130_fd_sc_hd__buf_1 _13929_ (.A(_10845_),
    .X(_11065_));
 sky130_fd_sc_hd__o221a_2 _13930_ (.A1(eoi[11]),
    .A2(_11059_),
    .B1(_11060_),
    .B2(_11064_),
    .C1(_11065_),
    .X(_03844_));
 sky130_fd_sc_hd__nor3_2 _13931_ (.A(\irq_mask[10] ),
    .B(_10550_),
    .C(_11050_),
    .Y(_11066_));
 sky130_fd_sc_hd__o221a_2 _13932_ (.A1(eoi[10]),
    .A2(_11059_),
    .B1(_11060_),
    .B2(_11066_),
    .C1(_11065_),
    .X(_03843_));
 sky130_fd_sc_hd__and3_2 _13933_ (.A(_10547_),
    .B(\irq_pending[9] ),
    .C(_11063_),
    .X(_11067_));
 sky130_fd_sc_hd__o221a_2 _13934_ (.A1(eoi[9]),
    .A2(_11059_),
    .B1(_11060_),
    .B2(_11067_),
    .C1(_11065_),
    .X(_03842_));
 sky130_fd_sc_hd__nor3_2 _13935_ (.A(\irq_mask[8] ),
    .B(_10549_),
    .C(_11027_),
    .Y(_11068_));
 sky130_fd_sc_hd__o221a_2 _13936_ (.A1(eoi[8]),
    .A2(_11059_),
    .B1(_11060_),
    .B2(_11068_),
    .C1(_11065_),
    .X(_03841_));
 sky130_fd_sc_hd__buf_1 _13937_ (.A(_11021_),
    .X(_11069_));
 sky130_fd_sc_hd__buf_1 _13938_ (.A(_11024_),
    .X(_11070_));
 sky130_fd_sc_hd__and3_2 _13939_ (.A(_10529_),
    .B(\irq_pending[7] ),
    .C(_11063_),
    .X(_11071_));
 sky130_fd_sc_hd__o221a_2 _13940_ (.A1(eoi[7]),
    .A2(_11069_),
    .B1(_11070_),
    .B2(_11071_),
    .C1(_11065_),
    .X(_03840_));
 sky130_fd_sc_hd__nor3_2 _13941_ (.A(\irq_mask[6] ),
    .B(_10531_),
    .C(_11027_),
    .Y(_11072_));
 sky130_fd_sc_hd__o221a_2 _13942_ (.A1(eoi[6]),
    .A2(_11069_),
    .B1(_11070_),
    .B2(_11072_),
    .C1(_11065_),
    .X(_03839_));
 sky130_fd_sc_hd__and3_2 _13943_ (.A(_10528_),
    .B(\irq_pending[5] ),
    .C(_11063_),
    .X(_11073_));
 sky130_fd_sc_hd__buf_1 _13944_ (.A(_10845_),
    .X(_11074_));
 sky130_fd_sc_hd__o221a_2 _13945_ (.A1(eoi[5]),
    .A2(_11069_),
    .B1(_11070_),
    .B2(_11073_),
    .C1(_11074_),
    .X(_03838_));
 sky130_fd_sc_hd__nor3_2 _13946_ (.A(\irq_mask[4] ),
    .B(_10530_),
    .C(_11027_),
    .Y(_11075_));
 sky130_fd_sc_hd__o221a_2 _13947_ (.A1(eoi[4]),
    .A2(_11069_),
    .B1(_11070_),
    .B2(_11075_),
    .C1(_11074_),
    .X(_03837_));
 sky130_fd_sc_hd__nor3_2 _13948_ (.A(\irq_mask[3] ),
    .B(_10513_),
    .C(_11027_),
    .Y(_11076_));
 sky130_fd_sc_hd__o221a_2 _13949_ (.A1(eoi[3]),
    .A2(_11069_),
    .B1(_11070_),
    .B2(_11076_),
    .C1(_11074_),
    .X(_03836_));
 sky130_fd_sc_hd__and3_2 _13950_ (.A(_10511_),
    .B(\irq_pending[2] ),
    .C(_11063_),
    .X(_11077_));
 sky130_fd_sc_hd__o221a_2 _13951_ (.A1(eoi[2]),
    .A2(_11069_),
    .B1(_11070_),
    .B2(_11077_),
    .C1(_11074_),
    .X(_03835_));
 sky130_fd_sc_hd__and3_2 _13952_ (.A(_10510_),
    .B(\irq_pending[1] ),
    .C(_11063_),
    .X(_11078_));
 sky130_fd_sc_hd__o221a_2 _13953_ (.A1(eoi[1]),
    .A2(_11022_),
    .B1(_11025_),
    .B2(_11078_),
    .C1(_11074_),
    .X(_03834_));
 sky130_vsdinv _13954_ (.A(\irq_mask[0] ),
    .Y(_11079_));
 sky130_fd_sc_hd__buf_1 _13955_ (.A(_10469_),
    .X(_11080_));
 sky130_fd_sc_hd__and3_2 _13956_ (.A(_11079_),
    .B(\irq_pending[0] ),
    .C(_11080_),
    .X(_11081_));
 sky130_fd_sc_hd__o221a_2 _13957_ (.A1(eoi[0]),
    .A2(_11022_),
    .B1(_11025_),
    .B2(_11081_),
    .C1(_11074_),
    .X(_03833_));
 sky130_vsdinv _13958_ (.A(_10639_),
    .Y(_11082_));
 sky130_fd_sc_hd__or2_2 _13959_ (.A(_11082_),
    .B(_10638_),
    .X(_11083_));
 sky130_fd_sc_hd__buf_1 _13960_ (.A(_10639_),
    .X(_11084_));
 sky130_fd_sc_hd__buf_1 _13961_ (.A(_11084_),
    .X(_11085_));
 sky130_fd_sc_hd__nor2_2 _13962_ (.A(instr_ecall_ebreak),
    .B(pcpi_timeout),
    .Y(_00311_));
 sky130_fd_sc_hd__nand2_2 _13963_ (.A(_10623_),
    .B(_00311_),
    .Y(_11086_));
 sky130_fd_sc_hd__a31o_2 _13964_ (.A1(_11085_),
    .A2(_00310_),
    .A3(_11086_),
    .B1(_10774_),
    .X(_11087_));
 sky130_fd_sc_hd__a21oi_2 _13965_ (.A1(_10569_),
    .A2(_11083_),
    .B1(_11087_),
    .Y(_03832_));
 sky130_fd_sc_hd__inv_2 _13966_ (.A(_10452_),
    .Y(_00290_));
 sky130_fd_sc_hd__o31a_2 _13967_ (.A1(mem_do_wdata),
    .A2(_10484_),
    .A3(mem_valid),
    .B1(_00290_),
    .X(_11088_));
 sky130_fd_sc_hd__a21oi_2 _13968_ (.A1(mem_valid),
    .A2(_10450_),
    .B1(_11088_),
    .Y(_11089_));
 sky130_vsdinv _13969_ (.A(mem_valid),
    .Y(_11090_));
 sky130_fd_sc_hd__o22a_2 _13970_ (.A1(trap),
    .A2(_11089_),
    .B1(_11090_),
    .B2(mem_ready),
    .X(_11091_));
 sky130_fd_sc_hd__nor2_2 _13971_ (.A(_10791_),
    .B(_11091_),
    .Y(_03831_));
 sky130_fd_sc_hd__or4_2 _13972_ (.A(\irq_pending[21] ),
    .B(\irq_pending[20] ),
    .C(\irq_pending[23] ),
    .D(\irq_pending[22] ),
    .X(_11092_));
 sky130_fd_sc_hd__or4_2 _13973_ (.A(\irq_pending[17] ),
    .B(\irq_pending[16] ),
    .C(\irq_pending[19] ),
    .D(\irq_pending[18] ),
    .X(_11093_));
 sky130_fd_sc_hd__or4_2 _13974_ (.A(\irq_pending[29] ),
    .B(\irq_pending[28] ),
    .C(\irq_pending[31] ),
    .D(\irq_pending[30] ),
    .X(_11094_));
 sky130_fd_sc_hd__or4_2 _13975_ (.A(\irq_pending[25] ),
    .B(\irq_pending[24] ),
    .C(\irq_pending[27] ),
    .D(\irq_pending[26] ),
    .X(_11095_));
 sky130_fd_sc_hd__or4_2 _13976_ (.A(_11092_),
    .B(_11093_),
    .C(_11094_),
    .D(_11095_),
    .X(_11096_));
 sky130_fd_sc_hd__or4_2 _13977_ (.A(\irq_pending[5] ),
    .B(\irq_pending[4] ),
    .C(\irq_pending[7] ),
    .D(\irq_pending[6] ),
    .X(_11097_));
 sky130_fd_sc_hd__or4_2 _13978_ (.A(\irq_pending[1] ),
    .B(\irq_pending[0] ),
    .C(\irq_pending[3] ),
    .D(\irq_pending[2] ),
    .X(_11098_));
 sky130_fd_sc_hd__or4_2 _13979_ (.A(\irq_pending[13] ),
    .B(\irq_pending[12] ),
    .C(\irq_pending[15] ),
    .D(\irq_pending[14] ),
    .X(_11099_));
 sky130_fd_sc_hd__or4_2 _13980_ (.A(\irq_pending[9] ),
    .B(\irq_pending[8] ),
    .C(\irq_pending[11] ),
    .D(\irq_pending[10] ),
    .X(_11100_));
 sky130_fd_sc_hd__or4_2 _13981_ (.A(_11097_),
    .B(_11098_),
    .C(_11099_),
    .D(_11100_),
    .X(_11101_));
 sky130_fd_sc_hd__or2_2 _13982_ (.A(_11096_),
    .B(_11101_),
    .X(_11102_));
 sky130_fd_sc_hd__inv_2 _13983_ (.A(_11102_),
    .Y(_02410_));
 sky130_fd_sc_hd__buf_1 _13984_ (.A(_10563_),
    .X(_00308_));
 sky130_fd_sc_hd__or2_2 _13985_ (.A(_10475_),
    .B(_00308_),
    .X(_11103_));
 sky130_fd_sc_hd__or2_2 _13986_ (.A(_10564_),
    .B(_11103_),
    .X(_11104_));
 sky130_fd_sc_hd__nor3_2 _13987_ (.A(_00322_),
    .B(_11102_),
    .C(_11104_),
    .Y(_03830_));
 sky130_fd_sc_hd__or3_2 _13988_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(instr_sltu),
    .C(instr_slt),
    .X(_11105_));
 sky130_fd_sc_hd__buf_1 _13989_ (.A(_10463_),
    .X(_11106_));
 sky130_fd_sc_hd__buf_1 _13990_ (.A(_10760_),
    .X(_11107_));
 sky130_fd_sc_hd__o311a_2 _13991_ (.A1(instr_sltiu),
    .A2(instr_slti),
    .A3(_11105_),
    .B1(_11106_),
    .C1(_11107_),
    .X(_03829_));
 sky130_fd_sc_hd__inv_2 _13992_ (.A(_10671_),
    .Y(_00297_));
 sky130_fd_sc_hd__or2_2 _13993_ (.A(mem_do_prefetch),
    .B(_10454_),
    .X(_11108_));
 sky130_fd_sc_hd__or2_2 _13994_ (.A(_00297_),
    .B(_11108_),
    .X(_11109_));
 sky130_vsdinv _13995_ (.A(_11109_),
    .Y(_03828_));
 sky130_fd_sc_hd__nor2_2 _13996_ (.A(_11017_),
    .B(_10806_),
    .Y(_03827_));
 sky130_fd_sc_hd__buf_1 _13997_ (.A(_10444_),
    .X(_11110_));
 sky130_fd_sc_hd__buf_1 _13998_ (.A(_11110_),
    .X(_11111_));
 sky130_fd_sc_hd__and2_2 _13999_ (.A(_11111_),
    .B(_02435_),
    .X(_03826_));
 sky130_fd_sc_hd__and2_2 _14000_ (.A(_11111_),
    .B(_02434_),
    .X(_03825_));
 sky130_fd_sc_hd__and2_2 _14001_ (.A(_11111_),
    .B(_02432_),
    .X(_03824_));
 sky130_fd_sc_hd__and2_2 _14002_ (.A(_11111_),
    .B(_02431_),
    .X(_03823_));
 sky130_fd_sc_hd__and2_2 _14003_ (.A(_11111_),
    .B(_02430_),
    .X(_03822_));
 sky130_fd_sc_hd__buf_1 _14004_ (.A(_11110_),
    .X(_11112_));
 sky130_fd_sc_hd__and2_2 _14005_ (.A(_11112_),
    .B(_02429_),
    .X(_03821_));
 sky130_fd_sc_hd__and2_2 _14006_ (.A(_11112_),
    .B(_02428_),
    .X(_03820_));
 sky130_fd_sc_hd__and2_2 _14007_ (.A(_11112_),
    .B(_02427_),
    .X(_03819_));
 sky130_fd_sc_hd__and2_2 _14008_ (.A(_11112_),
    .B(_02426_),
    .X(_03818_));
 sky130_fd_sc_hd__and2_2 _14009_ (.A(_11112_),
    .B(_02425_),
    .X(_03817_));
 sky130_fd_sc_hd__and2_2 _14010_ (.A(_11112_),
    .B(_02424_),
    .X(_03816_));
 sky130_fd_sc_hd__buf_1 _14011_ (.A(_11110_),
    .X(_11113_));
 sky130_fd_sc_hd__and2_2 _14012_ (.A(_11113_),
    .B(_02423_),
    .X(_03815_));
 sky130_fd_sc_hd__and2_2 _14013_ (.A(_11113_),
    .B(_02421_),
    .X(_03814_));
 sky130_fd_sc_hd__and2_2 _14014_ (.A(_11113_),
    .B(_02420_),
    .X(_03813_));
 sky130_fd_sc_hd__and2_2 _14015_ (.A(_11113_),
    .B(_02419_),
    .X(_03812_));
 sky130_fd_sc_hd__and2_2 _14016_ (.A(_11113_),
    .B(_02418_),
    .X(_03811_));
 sky130_fd_sc_hd__and2_2 _14017_ (.A(_11113_),
    .B(_02417_),
    .X(_03810_));
 sky130_fd_sc_hd__buf_1 _14018_ (.A(_10444_),
    .X(_11114_));
 sky130_fd_sc_hd__buf_1 _14019_ (.A(_11114_),
    .X(_11115_));
 sky130_fd_sc_hd__and2_2 _14020_ (.A(_11115_),
    .B(_02416_),
    .X(_03809_));
 sky130_fd_sc_hd__and2_2 _14021_ (.A(_11115_),
    .B(_02415_),
    .X(_03808_));
 sky130_fd_sc_hd__and2_2 _14022_ (.A(_11115_),
    .B(_02414_),
    .X(_03807_));
 sky130_fd_sc_hd__and2_2 _14023_ (.A(_11115_),
    .B(_02413_),
    .X(_03806_));
 sky130_fd_sc_hd__and2_2 _14024_ (.A(_11115_),
    .B(_02412_),
    .X(_03805_));
 sky130_fd_sc_hd__and2_2 _14025_ (.A(_11115_),
    .B(_02442_),
    .X(_03804_));
 sky130_fd_sc_hd__buf_1 _14026_ (.A(_11114_),
    .X(_11116_));
 sky130_fd_sc_hd__and2_2 _14027_ (.A(_11116_),
    .B(_02441_),
    .X(_03803_));
 sky130_fd_sc_hd__and2_2 _14028_ (.A(_11116_),
    .B(_02440_),
    .X(_03802_));
 sky130_fd_sc_hd__and2_2 _14029_ (.A(_11116_),
    .B(_02439_),
    .X(_03801_));
 sky130_fd_sc_hd__and2_2 _14030_ (.A(_11116_),
    .B(_02438_),
    .X(_03800_));
 sky130_fd_sc_hd__and2_2 _14031_ (.A(_11116_),
    .B(_02437_),
    .X(_03799_));
 sky130_fd_sc_hd__and2_2 _14032_ (.A(_11116_),
    .B(_02436_),
    .X(_03798_));
 sky130_fd_sc_hd__buf_1 _14033_ (.A(_11114_),
    .X(_11117_));
 sky130_fd_sc_hd__and2_2 _14034_ (.A(_11117_),
    .B(_02433_),
    .X(_03797_));
 sky130_fd_sc_hd__and2_2 _14035_ (.A(_11117_),
    .B(_02422_),
    .X(_03796_));
 sky130_fd_sc_hd__and2_2 _14036_ (.A(_11117_),
    .B(_02411_),
    .X(_03795_));
 sky130_vsdinv _14037_ (.A(\count_cycle[62] ),
    .Y(_11118_));
 sky130_vsdinv _14038_ (.A(\count_cycle[61] ),
    .Y(_11119_));
 sky130_vsdinv _14039_ (.A(\count_cycle[60] ),
    .Y(_11120_));
 sky130_vsdinv _14040_ (.A(\count_cycle[59] ),
    .Y(_11121_));
 sky130_vsdinv _14041_ (.A(\count_cycle[58] ),
    .Y(_11122_));
 sky130_vsdinv _14042_ (.A(\count_cycle[57] ),
    .Y(_11123_));
 sky130_vsdinv _14043_ (.A(\count_cycle[56] ),
    .Y(_11124_));
 sky130_vsdinv _14044_ (.A(\count_cycle[55] ),
    .Y(_11125_));
 sky130_vsdinv _14045_ (.A(\count_cycle[54] ),
    .Y(_11126_));
 sky130_vsdinv _14046_ (.A(\count_cycle[53] ),
    .Y(_11127_));
 sky130_vsdinv _14047_ (.A(\count_cycle[52] ),
    .Y(_11128_));
 sky130_vsdinv _14048_ (.A(\count_cycle[51] ),
    .Y(_11129_));
 sky130_vsdinv _14049_ (.A(\count_cycle[50] ),
    .Y(_11130_));
 sky130_vsdinv _14050_ (.A(\count_cycle[49] ),
    .Y(_11131_));
 sky130_vsdinv _14051_ (.A(\count_cycle[48] ),
    .Y(_11132_));
 sky130_vsdinv _14052_ (.A(\count_cycle[47] ),
    .Y(_11133_));
 sky130_vsdinv _14053_ (.A(\count_cycle[46] ),
    .Y(_11134_));
 sky130_vsdinv _14054_ (.A(\count_cycle[45] ),
    .Y(_11135_));
 sky130_vsdinv _14055_ (.A(\count_cycle[44] ),
    .Y(_11136_));
 sky130_vsdinv _14056_ (.A(\count_cycle[43] ),
    .Y(_11137_));
 sky130_vsdinv _14057_ (.A(\count_cycle[42] ),
    .Y(_11138_));
 sky130_vsdinv _14058_ (.A(\count_cycle[41] ),
    .Y(_11139_));
 sky130_vsdinv _14059_ (.A(\count_cycle[40] ),
    .Y(_11140_));
 sky130_vsdinv _14060_ (.A(\count_cycle[39] ),
    .Y(_11141_));
 sky130_vsdinv _14061_ (.A(\count_cycle[38] ),
    .Y(_11142_));
 sky130_vsdinv _14062_ (.A(\count_cycle[37] ),
    .Y(_11143_));
 sky130_vsdinv _14063_ (.A(\count_cycle[36] ),
    .Y(_11144_));
 sky130_vsdinv _14064_ (.A(\count_cycle[35] ),
    .Y(_11145_));
 sky130_vsdinv _14065_ (.A(\count_cycle[34] ),
    .Y(_11146_));
 sky130_vsdinv _14066_ (.A(\count_cycle[33] ),
    .Y(_11147_));
 sky130_vsdinv _14067_ (.A(\count_cycle[32] ),
    .Y(_11148_));
 sky130_vsdinv _14068_ (.A(\count_cycle[31] ),
    .Y(_02055_));
 sky130_fd_sc_hd__inv_2 _14069_ (.A(\count_cycle[30] ),
    .Y(_02046_));
 sky130_vsdinv _14070_ (.A(\count_cycle[29] ),
    .Y(_02037_));
 sky130_fd_sc_hd__inv_2 _14071_ (.A(\count_cycle[28] ),
    .Y(_02028_));
 sky130_vsdinv _14072_ (.A(\count_cycle[27] ),
    .Y(_02019_));
 sky130_fd_sc_hd__inv_2 _14073_ (.A(\count_cycle[26] ),
    .Y(_02010_));
 sky130_vsdinv _14074_ (.A(\count_cycle[25] ),
    .Y(_02001_));
 sky130_fd_sc_hd__inv_2 _14075_ (.A(\count_cycle[24] ),
    .Y(_01992_));
 sky130_vsdinv _14076_ (.A(\count_cycle[23] ),
    .Y(_01983_));
 sky130_fd_sc_hd__inv_2 _14077_ (.A(\count_cycle[22] ),
    .Y(_01974_));
 sky130_vsdinv _14078_ (.A(\count_cycle[21] ),
    .Y(_01965_));
 sky130_fd_sc_hd__inv_2 _14079_ (.A(\count_cycle[20] ),
    .Y(_01956_));
 sky130_vsdinv _14080_ (.A(\count_cycle[19] ),
    .Y(_01947_));
 sky130_fd_sc_hd__inv_2 _14081_ (.A(\count_cycle[18] ),
    .Y(_01938_));
 sky130_vsdinv _14082_ (.A(\count_cycle[17] ),
    .Y(_01929_));
 sky130_fd_sc_hd__inv_2 _14083_ (.A(\count_cycle[16] ),
    .Y(_01920_));
 sky130_vsdinv _14084_ (.A(\count_cycle[15] ),
    .Y(_01911_));
 sky130_fd_sc_hd__inv_2 _14085_ (.A(\count_cycle[14] ),
    .Y(_01898_));
 sky130_vsdinv _14086_ (.A(\count_cycle[13] ),
    .Y(_01885_));
 sky130_fd_sc_hd__inv_2 _14087_ (.A(\count_cycle[12] ),
    .Y(_01872_));
 sky130_vsdinv _14088_ (.A(\count_cycle[11] ),
    .Y(_01859_));
 sky130_fd_sc_hd__inv_2 _14089_ (.A(\count_cycle[10] ),
    .Y(_01846_));
 sky130_vsdinv _14090_ (.A(\count_cycle[9] ),
    .Y(_01833_));
 sky130_fd_sc_hd__inv_2 _14091_ (.A(\count_cycle[8] ),
    .Y(_01820_));
 sky130_vsdinv _14092_ (.A(\count_cycle[7] ),
    .Y(_01806_));
 sky130_fd_sc_hd__inv_2 _14093_ (.A(\count_cycle[6] ),
    .Y(_01793_));
 sky130_vsdinv _14094_ (.A(\count_cycle[5] ),
    .Y(_01780_));
 sky130_vsdinv _14095_ (.A(\count_cycle[4] ),
    .Y(_01767_));
 sky130_fd_sc_hd__inv_2 _14096_ (.A(\count_cycle[0] ),
    .Y(_02559_));
 sky130_fd_sc_hd__inv_2 _14097_ (.A(\count_cycle[1] ),
    .Y(_01728_));
 sky130_fd_sc_hd__inv_2 _14098_ (.A(\count_cycle[2] ),
    .Y(_01741_));
 sky130_fd_sc_hd__inv_2 _14099_ (.A(\count_cycle[3] ),
    .Y(_01754_));
 sky130_fd_sc_hd__or4_2 _14100_ (.A(_02559_),
    .B(_01728_),
    .C(_01741_),
    .D(_01754_),
    .X(_11149_));
 sky130_fd_sc_hd__or2_2 _14101_ (.A(_01767_),
    .B(_11149_),
    .X(_11150_));
 sky130_fd_sc_hd__or2_2 _14102_ (.A(_01780_),
    .B(_11150_),
    .X(_11151_));
 sky130_fd_sc_hd__or2_2 _14103_ (.A(_01793_),
    .B(_11151_),
    .X(_11152_));
 sky130_fd_sc_hd__or2_2 _14104_ (.A(_01806_),
    .B(_11152_),
    .X(_11153_));
 sky130_fd_sc_hd__or2_2 _14105_ (.A(_01820_),
    .B(_11153_),
    .X(_11154_));
 sky130_fd_sc_hd__or2_2 _14106_ (.A(_01833_),
    .B(_11154_),
    .X(_11155_));
 sky130_fd_sc_hd__or2_2 _14107_ (.A(_01846_),
    .B(_11155_),
    .X(_11156_));
 sky130_fd_sc_hd__or2_2 _14108_ (.A(_01859_),
    .B(_11156_),
    .X(_11157_));
 sky130_fd_sc_hd__or2_2 _14109_ (.A(_01872_),
    .B(_11157_),
    .X(_11158_));
 sky130_fd_sc_hd__or2_2 _14110_ (.A(_01885_),
    .B(_11158_),
    .X(_11159_));
 sky130_fd_sc_hd__or2_2 _14111_ (.A(_01898_),
    .B(_11159_),
    .X(_11160_));
 sky130_fd_sc_hd__or2_2 _14112_ (.A(_01911_),
    .B(_11160_),
    .X(_11161_));
 sky130_fd_sc_hd__or2_2 _14113_ (.A(_01920_),
    .B(_11161_),
    .X(_11162_));
 sky130_fd_sc_hd__or2_2 _14114_ (.A(_01929_),
    .B(_11162_),
    .X(_11163_));
 sky130_fd_sc_hd__or2_2 _14115_ (.A(_01938_),
    .B(_11163_),
    .X(_11164_));
 sky130_fd_sc_hd__or2_2 _14116_ (.A(_01947_),
    .B(_11164_),
    .X(_11165_));
 sky130_fd_sc_hd__or2_2 _14117_ (.A(_01956_),
    .B(_11165_),
    .X(_11166_));
 sky130_fd_sc_hd__or2_2 _14118_ (.A(_01965_),
    .B(_11166_),
    .X(_11167_));
 sky130_fd_sc_hd__or2_2 _14119_ (.A(_01974_),
    .B(_11167_),
    .X(_11168_));
 sky130_fd_sc_hd__or2_2 _14120_ (.A(_01983_),
    .B(_11168_),
    .X(_11169_));
 sky130_fd_sc_hd__or2_2 _14121_ (.A(_01992_),
    .B(_11169_),
    .X(_11170_));
 sky130_fd_sc_hd__or2_2 _14122_ (.A(_02001_),
    .B(_11170_),
    .X(_11171_));
 sky130_fd_sc_hd__or2_2 _14123_ (.A(_02010_),
    .B(_11171_),
    .X(_11172_));
 sky130_fd_sc_hd__or2_2 _14124_ (.A(_02019_),
    .B(_11172_),
    .X(_11173_));
 sky130_fd_sc_hd__or2_2 _14125_ (.A(_02028_),
    .B(_11173_),
    .X(_11174_));
 sky130_fd_sc_hd__or2_2 _14126_ (.A(_02037_),
    .B(_11174_),
    .X(_11175_));
 sky130_fd_sc_hd__or2_2 _14127_ (.A(_02046_),
    .B(_11175_),
    .X(_11176_));
 sky130_fd_sc_hd__or2_2 _14128_ (.A(_02055_),
    .B(_11176_),
    .X(_11177_));
 sky130_fd_sc_hd__or2_2 _14129_ (.A(_11148_),
    .B(_11177_),
    .X(_11178_));
 sky130_fd_sc_hd__or2_2 _14130_ (.A(_11147_),
    .B(_11178_),
    .X(_11179_));
 sky130_fd_sc_hd__or2_2 _14131_ (.A(_11146_),
    .B(_11179_),
    .X(_11180_));
 sky130_fd_sc_hd__or2_2 _14132_ (.A(_11145_),
    .B(_11180_),
    .X(_11181_));
 sky130_fd_sc_hd__or2_2 _14133_ (.A(_11144_),
    .B(_11181_),
    .X(_11182_));
 sky130_fd_sc_hd__or2_2 _14134_ (.A(_11143_),
    .B(_11182_),
    .X(_11183_));
 sky130_fd_sc_hd__or2_2 _14135_ (.A(_11142_),
    .B(_11183_),
    .X(_11184_));
 sky130_fd_sc_hd__or2_2 _14136_ (.A(_11141_),
    .B(_11184_),
    .X(_11185_));
 sky130_fd_sc_hd__or2_2 _14137_ (.A(_11140_),
    .B(_11185_),
    .X(_11186_));
 sky130_fd_sc_hd__or2_2 _14138_ (.A(_11139_),
    .B(_11186_),
    .X(_11187_));
 sky130_fd_sc_hd__or2_2 _14139_ (.A(_11138_),
    .B(_11187_),
    .X(_11188_));
 sky130_fd_sc_hd__or2_2 _14140_ (.A(_11137_),
    .B(_11188_),
    .X(_11189_));
 sky130_fd_sc_hd__or2_2 _14141_ (.A(_11136_),
    .B(_11189_),
    .X(_11190_));
 sky130_fd_sc_hd__or2_2 _14142_ (.A(_11135_),
    .B(_11190_),
    .X(_11191_));
 sky130_fd_sc_hd__or2_2 _14143_ (.A(_11134_),
    .B(_11191_),
    .X(_11192_));
 sky130_fd_sc_hd__or2_2 _14144_ (.A(_11133_),
    .B(_11192_),
    .X(_11193_));
 sky130_fd_sc_hd__or2_2 _14145_ (.A(_11132_),
    .B(_11193_),
    .X(_11194_));
 sky130_fd_sc_hd__or2_2 _14146_ (.A(_11131_),
    .B(_11194_),
    .X(_11195_));
 sky130_fd_sc_hd__or2_2 _14147_ (.A(_11130_),
    .B(_11195_),
    .X(_11196_));
 sky130_fd_sc_hd__or2_2 _14148_ (.A(_11129_),
    .B(_11196_),
    .X(_11197_));
 sky130_fd_sc_hd__or2_2 _14149_ (.A(_11128_),
    .B(_11197_),
    .X(_11198_));
 sky130_fd_sc_hd__or2_2 _14150_ (.A(_11127_),
    .B(_11198_),
    .X(_11199_));
 sky130_fd_sc_hd__or2_2 _14151_ (.A(_11126_),
    .B(_11199_),
    .X(_11200_));
 sky130_fd_sc_hd__or2_2 _14152_ (.A(_11125_),
    .B(_11200_),
    .X(_11201_));
 sky130_fd_sc_hd__or2_2 _14153_ (.A(_11124_),
    .B(_11201_),
    .X(_11202_));
 sky130_fd_sc_hd__or2_2 _14154_ (.A(_11123_),
    .B(_11202_),
    .X(_11203_));
 sky130_fd_sc_hd__or2_2 _14155_ (.A(_11122_),
    .B(_11203_),
    .X(_11204_));
 sky130_fd_sc_hd__or2_2 _14156_ (.A(_11121_),
    .B(_11204_),
    .X(_11205_));
 sky130_fd_sc_hd__or2_2 _14157_ (.A(_11120_),
    .B(_11205_),
    .X(_11206_));
 sky130_fd_sc_hd__or2_2 _14158_ (.A(_11119_),
    .B(_11206_),
    .X(_11207_));
 sky130_fd_sc_hd__or2_2 _14159_ (.A(_11118_),
    .B(_11207_),
    .X(_11208_));
 sky130_vsdinv _14160_ (.A(_11208_),
    .Y(_11209_));
 sky130_vsdinv _14161_ (.A(\count_cycle[63] ),
    .Y(_11210_));
 sky130_fd_sc_hd__o221a_2 _14162_ (.A1(\count_cycle[63] ),
    .A2(_11209_),
    .B1(_11210_),
    .B2(_11208_),
    .C1(_11106_),
    .X(_03794_));
 sky130_fd_sc_hd__a211oi_2 _14163_ (.A1(_11118_),
    .A2(_11207_),
    .B1(_11014_),
    .C1(_11209_),
    .Y(_03793_));
 sky130_vsdinv _14164_ (.A(_11206_),
    .Y(_11211_));
 sky130_fd_sc_hd__o211a_2 _14165_ (.A1(\count_cycle[61] ),
    .A2(_11211_),
    .B1(_11016_),
    .C1(_11207_),
    .X(_03792_));
 sky130_fd_sc_hd__a211oi_2 _14166_ (.A1(_11120_),
    .A2(_11205_),
    .B1(_11014_),
    .C1(_11211_),
    .Y(_03791_));
 sky130_vsdinv _14167_ (.A(_11204_),
    .Y(_11212_));
 sky130_fd_sc_hd__o211a_2 _14168_ (.A1(\count_cycle[59] ),
    .A2(_11212_),
    .B1(_11016_),
    .C1(_11205_),
    .X(_03790_));
 sky130_fd_sc_hd__a211oi_2 _14169_ (.A1(_11122_),
    .A2(_11203_),
    .B1(_11014_),
    .C1(_11212_),
    .Y(_03789_));
 sky130_vsdinv _14170_ (.A(_11202_),
    .Y(_11213_));
 sky130_fd_sc_hd__o211a_2 _14171_ (.A1(\count_cycle[57] ),
    .A2(_11213_),
    .B1(_11016_),
    .C1(_11203_),
    .X(_03788_));
 sky130_fd_sc_hd__a211oi_2 _14172_ (.A1(_11124_),
    .A2(_11201_),
    .B1(_11014_),
    .C1(_11213_),
    .Y(_03787_));
 sky130_vsdinv _14173_ (.A(_11200_),
    .Y(_11214_));
 sky130_fd_sc_hd__o211a_2 _14174_ (.A1(\count_cycle[55] ),
    .A2(_11214_),
    .B1(_11016_),
    .C1(_11201_),
    .X(_03786_));
 sky130_fd_sc_hd__a211oi_2 _14175_ (.A1(_11126_),
    .A2(_11199_),
    .B1(_11014_),
    .C1(_11214_),
    .Y(_03785_));
 sky130_vsdinv _14176_ (.A(_11198_),
    .Y(_11215_));
 sky130_fd_sc_hd__buf_1 _14177_ (.A(_11007_),
    .X(_11216_));
 sky130_fd_sc_hd__o211a_2 _14178_ (.A1(\count_cycle[53] ),
    .A2(_11215_),
    .B1(_11216_),
    .C1(_11199_),
    .X(_03784_));
 sky130_fd_sc_hd__buf_1 _14179_ (.A(_10996_),
    .X(_11217_));
 sky130_fd_sc_hd__a211oi_2 _14180_ (.A1(_11128_),
    .A2(_11197_),
    .B1(_11217_),
    .C1(_11215_),
    .Y(_03783_));
 sky130_vsdinv _14181_ (.A(_11196_),
    .Y(_11218_));
 sky130_fd_sc_hd__o211a_2 _14182_ (.A1(\count_cycle[51] ),
    .A2(_11218_),
    .B1(_11216_),
    .C1(_11197_),
    .X(_03782_));
 sky130_fd_sc_hd__a211oi_2 _14183_ (.A1(_11130_),
    .A2(_11195_),
    .B1(_11217_),
    .C1(_11218_),
    .Y(_03781_));
 sky130_vsdinv _14184_ (.A(_11194_),
    .Y(_11219_));
 sky130_fd_sc_hd__o211a_2 _14185_ (.A1(\count_cycle[49] ),
    .A2(_11219_),
    .B1(_11216_),
    .C1(_11195_),
    .X(_03780_));
 sky130_fd_sc_hd__a211oi_2 _14186_ (.A1(_11132_),
    .A2(_11193_),
    .B1(_11217_),
    .C1(_11219_),
    .Y(_03779_));
 sky130_vsdinv _14187_ (.A(_11192_),
    .Y(_11220_));
 sky130_fd_sc_hd__o211a_2 _14188_ (.A1(\count_cycle[47] ),
    .A2(_11220_),
    .B1(_11216_),
    .C1(_11193_),
    .X(_03778_));
 sky130_fd_sc_hd__a211oi_2 _14189_ (.A1(_11134_),
    .A2(_11191_),
    .B1(_11217_),
    .C1(_11220_),
    .Y(_03777_));
 sky130_vsdinv _14190_ (.A(_11190_),
    .Y(_11221_));
 sky130_fd_sc_hd__o211a_2 _14191_ (.A1(\count_cycle[45] ),
    .A2(_11221_),
    .B1(_11216_),
    .C1(_11191_),
    .X(_03776_));
 sky130_fd_sc_hd__a211oi_2 _14192_ (.A1(_11136_),
    .A2(_11189_),
    .B1(_11217_),
    .C1(_11221_),
    .Y(_03775_));
 sky130_vsdinv _14193_ (.A(_11188_),
    .Y(_11222_));
 sky130_fd_sc_hd__o211a_2 _14194_ (.A1(\count_cycle[43] ),
    .A2(_11222_),
    .B1(_11216_),
    .C1(_11189_),
    .X(_03774_));
 sky130_fd_sc_hd__a211oi_2 _14195_ (.A1(_11138_),
    .A2(_11187_),
    .B1(_11217_),
    .C1(_11222_),
    .Y(_03773_));
 sky130_vsdinv _14196_ (.A(_11186_),
    .Y(_11223_));
 sky130_fd_sc_hd__buf_1 _14197_ (.A(_11007_),
    .X(_11224_));
 sky130_fd_sc_hd__o211a_2 _14198_ (.A1(\count_cycle[41] ),
    .A2(_11223_),
    .B1(_11224_),
    .C1(_11187_),
    .X(_03772_));
 sky130_fd_sc_hd__buf_1 _14199_ (.A(_10996_),
    .X(_11225_));
 sky130_fd_sc_hd__a211oi_2 _14200_ (.A1(_11140_),
    .A2(_11185_),
    .B1(_11225_),
    .C1(_11223_),
    .Y(_03771_));
 sky130_vsdinv _14201_ (.A(_11184_),
    .Y(_11226_));
 sky130_fd_sc_hd__o211a_2 _14202_ (.A1(\count_cycle[39] ),
    .A2(_11226_),
    .B1(_11224_),
    .C1(_11185_),
    .X(_03770_));
 sky130_fd_sc_hd__a211oi_2 _14203_ (.A1(_11142_),
    .A2(_11183_),
    .B1(_11225_),
    .C1(_11226_),
    .Y(_03769_));
 sky130_vsdinv _14204_ (.A(_11182_),
    .Y(_11227_));
 sky130_fd_sc_hd__o211a_2 _14205_ (.A1(\count_cycle[37] ),
    .A2(_11227_),
    .B1(_11224_),
    .C1(_11183_),
    .X(_03768_));
 sky130_fd_sc_hd__a211oi_2 _14206_ (.A1(_11144_),
    .A2(_11181_),
    .B1(_11225_),
    .C1(_11227_),
    .Y(_03767_));
 sky130_vsdinv _14207_ (.A(_11180_),
    .Y(_11228_));
 sky130_fd_sc_hd__o211a_2 _14208_ (.A1(\count_cycle[35] ),
    .A2(_11228_),
    .B1(_11224_),
    .C1(_11181_),
    .X(_03766_));
 sky130_fd_sc_hd__a211oi_2 _14209_ (.A1(_11146_),
    .A2(_11179_),
    .B1(_11225_),
    .C1(_11228_),
    .Y(_03765_));
 sky130_vsdinv _14210_ (.A(_11178_),
    .Y(_11229_));
 sky130_fd_sc_hd__o211a_2 _14211_ (.A1(\count_cycle[33] ),
    .A2(_11229_),
    .B1(_11224_),
    .C1(_11179_),
    .X(_03764_));
 sky130_fd_sc_hd__a211oi_2 _14212_ (.A1(_11148_),
    .A2(_11177_),
    .B1(_11225_),
    .C1(_11229_),
    .Y(_03763_));
 sky130_vsdinv _14213_ (.A(_11176_),
    .Y(_11230_));
 sky130_fd_sc_hd__o211a_2 _14214_ (.A1(\count_cycle[31] ),
    .A2(_11230_),
    .B1(_11224_),
    .C1(_11177_),
    .X(_03762_));
 sky130_fd_sc_hd__a211oi_2 _14215_ (.A1(_02046_),
    .A2(_11175_),
    .B1(_11225_),
    .C1(_11230_),
    .Y(_03761_));
 sky130_vsdinv _14216_ (.A(_11174_),
    .Y(_11231_));
 sky130_fd_sc_hd__buf_1 _14217_ (.A(_11007_),
    .X(_11232_));
 sky130_fd_sc_hd__o211a_2 _14218_ (.A1(\count_cycle[29] ),
    .A2(_11231_),
    .B1(_11232_),
    .C1(_11175_),
    .X(_03760_));
 sky130_fd_sc_hd__buf_1 _14219_ (.A(_10996_),
    .X(_11233_));
 sky130_fd_sc_hd__a211oi_2 _14220_ (.A1(_02028_),
    .A2(_11173_),
    .B1(_11233_),
    .C1(_11231_),
    .Y(_03759_));
 sky130_vsdinv _14221_ (.A(_11172_),
    .Y(_11234_));
 sky130_fd_sc_hd__o211a_2 _14222_ (.A1(\count_cycle[27] ),
    .A2(_11234_),
    .B1(_11232_),
    .C1(_11173_),
    .X(_03758_));
 sky130_fd_sc_hd__a211oi_2 _14223_ (.A1(_02010_),
    .A2(_11171_),
    .B1(_11233_),
    .C1(_11234_),
    .Y(_03757_));
 sky130_vsdinv _14224_ (.A(_11170_),
    .Y(_11235_));
 sky130_fd_sc_hd__o211a_2 _14225_ (.A1(\count_cycle[25] ),
    .A2(_11235_),
    .B1(_11232_),
    .C1(_11171_),
    .X(_03756_));
 sky130_fd_sc_hd__a211oi_2 _14226_ (.A1(_01992_),
    .A2(_11169_),
    .B1(_11233_),
    .C1(_11235_),
    .Y(_03755_));
 sky130_vsdinv _14227_ (.A(_11168_),
    .Y(_11236_));
 sky130_fd_sc_hd__o211a_2 _14228_ (.A1(\count_cycle[23] ),
    .A2(_11236_),
    .B1(_11232_),
    .C1(_11169_),
    .X(_03754_));
 sky130_fd_sc_hd__a211oi_2 _14229_ (.A1(_01974_),
    .A2(_11167_),
    .B1(_11233_),
    .C1(_11236_),
    .Y(_03753_));
 sky130_vsdinv _14230_ (.A(_11166_),
    .Y(_11237_));
 sky130_fd_sc_hd__o211a_2 _14231_ (.A1(\count_cycle[21] ),
    .A2(_11237_),
    .B1(_11232_),
    .C1(_11167_),
    .X(_03752_));
 sky130_fd_sc_hd__a211oi_2 _14232_ (.A1(_01956_),
    .A2(_11165_),
    .B1(_11233_),
    .C1(_11237_),
    .Y(_03751_));
 sky130_vsdinv _14233_ (.A(_11164_),
    .Y(_11238_));
 sky130_fd_sc_hd__o211a_2 _14234_ (.A1(\count_cycle[19] ),
    .A2(_11238_),
    .B1(_11232_),
    .C1(_11165_),
    .X(_03750_));
 sky130_fd_sc_hd__a211oi_2 _14235_ (.A1(_01938_),
    .A2(_11163_),
    .B1(_11233_),
    .C1(_11238_),
    .Y(_03749_));
 sky130_vsdinv _14236_ (.A(_11162_),
    .Y(_11239_));
 sky130_fd_sc_hd__buf_1 _14237_ (.A(_11007_),
    .X(_11240_));
 sky130_fd_sc_hd__o211a_2 _14238_ (.A1(\count_cycle[17] ),
    .A2(_11239_),
    .B1(_11240_),
    .C1(_11163_),
    .X(_03748_));
 sky130_fd_sc_hd__buf_1 _14239_ (.A(_10688_),
    .X(_11241_));
 sky130_fd_sc_hd__a211oi_2 _14240_ (.A1(_01920_),
    .A2(_11161_),
    .B1(_11241_),
    .C1(_11239_),
    .Y(_03747_));
 sky130_vsdinv _14241_ (.A(_11160_),
    .Y(_11242_));
 sky130_fd_sc_hd__o211a_2 _14242_ (.A1(\count_cycle[15] ),
    .A2(_11242_),
    .B1(_11240_),
    .C1(_11161_),
    .X(_03746_));
 sky130_fd_sc_hd__a211oi_2 _14243_ (.A1(_01898_),
    .A2(_11159_),
    .B1(_11241_),
    .C1(_11242_),
    .Y(_03745_));
 sky130_vsdinv _14244_ (.A(_11158_),
    .Y(_11243_));
 sky130_fd_sc_hd__o211a_2 _14245_ (.A1(\count_cycle[13] ),
    .A2(_11243_),
    .B1(_11240_),
    .C1(_11159_),
    .X(_03744_));
 sky130_fd_sc_hd__a211oi_2 _14246_ (.A1(_01872_),
    .A2(_11157_),
    .B1(_11241_),
    .C1(_11243_),
    .Y(_03743_));
 sky130_vsdinv _14247_ (.A(_11156_),
    .Y(_11244_));
 sky130_fd_sc_hd__o211a_2 _14248_ (.A1(\count_cycle[11] ),
    .A2(_11244_),
    .B1(_11240_),
    .C1(_11157_),
    .X(_03742_));
 sky130_fd_sc_hd__a211oi_2 _14249_ (.A1(_01846_),
    .A2(_11155_),
    .B1(_11241_),
    .C1(_11244_),
    .Y(_03741_));
 sky130_vsdinv _14250_ (.A(_11154_),
    .Y(_11245_));
 sky130_fd_sc_hd__o211a_2 _14251_ (.A1(\count_cycle[9] ),
    .A2(_11245_),
    .B1(_11240_),
    .C1(_11155_),
    .X(_03740_));
 sky130_fd_sc_hd__a211oi_2 _14252_ (.A1(_01820_),
    .A2(_11153_),
    .B1(_11241_),
    .C1(_11245_),
    .Y(_03739_));
 sky130_vsdinv _14253_ (.A(_11152_),
    .Y(_11246_));
 sky130_fd_sc_hd__o211a_2 _14254_ (.A1(\count_cycle[7] ),
    .A2(_11246_),
    .B1(_11240_),
    .C1(_11153_),
    .X(_03738_));
 sky130_fd_sc_hd__a211oi_2 _14255_ (.A1(_01793_),
    .A2(_11151_),
    .B1(_11241_),
    .C1(_11246_),
    .Y(_03737_));
 sky130_vsdinv _14256_ (.A(_11150_),
    .Y(_11247_));
 sky130_fd_sc_hd__o211a_2 _14257_ (.A1(\count_cycle[5] ),
    .A2(_11247_),
    .B1(_11110_),
    .C1(_11151_),
    .X(_03736_));
 sky130_vsdinv _14258_ (.A(_11149_),
    .Y(_11248_));
 sky130_fd_sc_hd__o211a_2 _14259_ (.A1(\count_cycle[4] ),
    .A2(_11248_),
    .B1(_11110_),
    .C1(_11150_),
    .X(_03735_));
 sky130_fd_sc_hd__o31a_2 _14260_ (.A1(_02559_),
    .A2(_01728_),
    .A3(_01741_),
    .B1(_01754_),
    .X(_11249_));
 sky130_fd_sc_hd__nor3_2 _14261_ (.A(_11017_),
    .B(_11248_),
    .C(_11249_),
    .Y(_03734_));
 sky130_fd_sc_hd__o21ai_2 _14262_ (.A1(_02559_),
    .A2(_01728_),
    .B1(_01741_),
    .Y(_11250_));
 sky130_fd_sc_hd__o311a_2 _14263_ (.A1(_02559_),
    .A2(_01728_),
    .A3(_01741_),
    .B1(_11106_),
    .C1(_11250_),
    .X(_03733_));
 sky130_fd_sc_hd__o221a_2 _14264_ (.A1(_02559_),
    .A2(_01728_),
    .B1(\count_cycle[0] ),
    .B2(\count_cycle[1] ),
    .C1(_11106_),
    .X(_03732_));
 sky130_fd_sc_hd__nor2_2 _14265_ (.A(_11017_),
    .B(\count_cycle[0] ),
    .Y(_03731_));
 sky130_vsdinv _14266_ (.A(\cpu_state[0] ),
    .Y(_11251_));
 sky130_fd_sc_hd__nor2_2 _14267_ (.A(_11017_),
    .B(_11251_),
    .Y(_03730_));
 sky130_fd_sc_hd__and2_2 _14268_ (.A(_11117_),
    .B(\pcpi_mul.active[0] ),
    .X(_03729_));
 sky130_fd_sc_hd__buf_1 _14269_ (.A(_10601_),
    .X(_03728_));
 sky130_fd_sc_hd__buf_1 _14270_ (.A(\latched_rd[3] ),
    .X(_11252_));
 sky130_vsdinv _14271_ (.A(\latched_rd[2] ),
    .Y(_11253_));
 sky130_fd_sc_hd__or3_2 _14272_ (.A(\latched_rd[4] ),
    .B(_11252_),
    .C(_11253_),
    .X(_11254_));
 sky130_vsdinv _14273_ (.A(latched_branch),
    .Y(_11255_));
 sky130_vsdinv _14274_ (.A(latched_store),
    .Y(_11256_));
 sky130_fd_sc_hd__and4_2 _14275_ (.A(_10649_),
    .B(_10648_),
    .C(_11255_),
    .D(_11256_),
    .X(_11257_));
 sky130_fd_sc_hd__or3_2 _14276_ (.A(\latched_rd[4] ),
    .B(\latched_rd[3] ),
    .C(\latched_rd[2] ),
    .X(_11258_));
 sky130_fd_sc_hd__nor3_2 _14277_ (.A(\latched_rd[0] ),
    .B(\latched_rd[1] ),
    .C(_11258_),
    .Y(_11259_));
 sky130_fd_sc_hd__or4_2 _14278_ (.A(_10474_),
    .B(_10508_),
    .C(_11257_),
    .D(_11259_),
    .X(_11260_));
 sky130_fd_sc_hd__or2b_2 _14279_ (.A(_11260_),
    .B_N(\latched_rd[1] ),
    .X(_11261_));
 sky130_fd_sc_hd__or2_2 _14280_ (.A(\latched_rd[0] ),
    .B(_11261_),
    .X(_11262_));
 sky130_fd_sc_hd__or2_2 _14281_ (.A(_11254_),
    .B(_11262_),
    .X(_11263_));
 sky130_fd_sc_hd__buf_1 _14282_ (.A(_11263_),
    .X(_11264_));
 sky130_fd_sc_hd__buf_1 _14283_ (.A(_11264_),
    .X(_11265_));
 sky130_fd_sc_hd__buf_1 _14284_ (.A(\cpuregs_wrdata[31] ),
    .X(_11266_));
 sky130_vsdinv _14285_ (.A(_11263_),
    .Y(_11267_));
 sky130_fd_sc_hd__buf_1 _14286_ (.A(_11267_),
    .X(_11268_));
 sky130_fd_sc_hd__buf_1 _14287_ (.A(_11268_),
    .X(_11269_));
 sky130_fd_sc_hd__a22o_2 _14288_ (.A1(\cpuregs[6][31] ),
    .A2(_11265_),
    .B1(_11266_),
    .B2(_11269_),
    .X(_03727_));
 sky130_fd_sc_hd__buf_1 _14289_ (.A(\cpuregs_wrdata[30] ),
    .X(_11270_));
 sky130_fd_sc_hd__a22o_2 _14290_ (.A1(\cpuregs[6][30] ),
    .A2(_11265_),
    .B1(_11270_),
    .B2(_11269_),
    .X(_03726_));
 sky130_fd_sc_hd__buf_1 _14291_ (.A(\cpuregs_wrdata[29] ),
    .X(_11271_));
 sky130_fd_sc_hd__a22o_2 _14292_ (.A1(\cpuregs[6][29] ),
    .A2(_11265_),
    .B1(_11271_),
    .B2(_11269_),
    .X(_03725_));
 sky130_fd_sc_hd__buf_1 _14293_ (.A(\cpuregs_wrdata[28] ),
    .X(_11272_));
 sky130_fd_sc_hd__a22o_2 _14294_ (.A1(\cpuregs[6][28] ),
    .A2(_11265_),
    .B1(_11272_),
    .B2(_11269_),
    .X(_03724_));
 sky130_fd_sc_hd__buf_1 _14295_ (.A(\cpuregs_wrdata[27] ),
    .X(_11273_));
 sky130_fd_sc_hd__a22o_2 _14296_ (.A1(\cpuregs[6][27] ),
    .A2(_11265_),
    .B1(_11273_),
    .B2(_11269_),
    .X(_03723_));
 sky130_fd_sc_hd__buf_1 _14297_ (.A(\cpuregs_wrdata[26] ),
    .X(_11274_));
 sky130_fd_sc_hd__a22o_2 _14298_ (.A1(\cpuregs[6][26] ),
    .A2(_11265_),
    .B1(_11274_),
    .B2(_11269_),
    .X(_03722_));
 sky130_fd_sc_hd__buf_1 _14299_ (.A(_11264_),
    .X(_11275_));
 sky130_fd_sc_hd__buf_1 _14300_ (.A(\cpuregs_wrdata[25] ),
    .X(_11276_));
 sky130_fd_sc_hd__buf_1 _14301_ (.A(_11268_),
    .X(_11277_));
 sky130_fd_sc_hd__a22o_2 _14302_ (.A1(\cpuregs[6][25] ),
    .A2(_11275_),
    .B1(_11276_),
    .B2(_11277_),
    .X(_03721_));
 sky130_fd_sc_hd__buf_1 _14303_ (.A(\cpuregs_wrdata[24] ),
    .X(_11278_));
 sky130_fd_sc_hd__a22o_2 _14304_ (.A1(\cpuregs[6][24] ),
    .A2(_11275_),
    .B1(_11278_),
    .B2(_11277_),
    .X(_03720_));
 sky130_fd_sc_hd__buf_1 _14305_ (.A(\cpuregs_wrdata[23] ),
    .X(_11279_));
 sky130_fd_sc_hd__a22o_2 _14306_ (.A1(\cpuregs[6][23] ),
    .A2(_11275_),
    .B1(_11279_),
    .B2(_11277_),
    .X(_03719_));
 sky130_fd_sc_hd__buf_1 _14307_ (.A(\cpuregs_wrdata[22] ),
    .X(_11280_));
 sky130_fd_sc_hd__a22o_2 _14308_ (.A1(\cpuregs[6][22] ),
    .A2(_11275_),
    .B1(_11280_),
    .B2(_11277_),
    .X(_03718_));
 sky130_fd_sc_hd__buf_1 _14309_ (.A(\cpuregs_wrdata[21] ),
    .X(_11281_));
 sky130_fd_sc_hd__a22o_2 _14310_ (.A1(\cpuregs[6][21] ),
    .A2(_11275_),
    .B1(_11281_),
    .B2(_11277_),
    .X(_03717_));
 sky130_fd_sc_hd__buf_1 _14311_ (.A(\cpuregs_wrdata[20] ),
    .X(_11282_));
 sky130_fd_sc_hd__a22o_2 _14312_ (.A1(\cpuregs[6][20] ),
    .A2(_11275_),
    .B1(_11282_),
    .B2(_11277_),
    .X(_03716_));
 sky130_fd_sc_hd__buf_1 _14313_ (.A(_11264_),
    .X(_11283_));
 sky130_fd_sc_hd__buf_1 _14314_ (.A(\cpuregs_wrdata[19] ),
    .X(_11284_));
 sky130_fd_sc_hd__buf_1 _14315_ (.A(_11268_),
    .X(_11285_));
 sky130_fd_sc_hd__a22o_2 _14316_ (.A1(\cpuregs[6][19] ),
    .A2(_11283_),
    .B1(_11284_),
    .B2(_11285_),
    .X(_03715_));
 sky130_fd_sc_hd__buf_1 _14317_ (.A(\cpuregs_wrdata[18] ),
    .X(_11286_));
 sky130_fd_sc_hd__a22o_2 _14318_ (.A1(\cpuregs[6][18] ),
    .A2(_11283_),
    .B1(_11286_),
    .B2(_11285_),
    .X(_03714_));
 sky130_fd_sc_hd__buf_1 _14319_ (.A(\cpuregs_wrdata[17] ),
    .X(_11287_));
 sky130_fd_sc_hd__a22o_2 _14320_ (.A1(\cpuregs[6][17] ),
    .A2(_11283_),
    .B1(_11287_),
    .B2(_11285_),
    .X(_03713_));
 sky130_fd_sc_hd__buf_1 _14321_ (.A(\cpuregs_wrdata[16] ),
    .X(_11288_));
 sky130_fd_sc_hd__a22o_2 _14322_ (.A1(\cpuregs[6][16] ),
    .A2(_11283_),
    .B1(_11288_),
    .B2(_11285_),
    .X(_03712_));
 sky130_fd_sc_hd__buf_1 _14323_ (.A(\cpuregs_wrdata[15] ),
    .X(_11289_));
 sky130_fd_sc_hd__a22o_2 _14324_ (.A1(\cpuregs[6][15] ),
    .A2(_11283_),
    .B1(_11289_),
    .B2(_11285_),
    .X(_03711_));
 sky130_fd_sc_hd__buf_1 _14325_ (.A(\cpuregs_wrdata[14] ),
    .X(_11290_));
 sky130_fd_sc_hd__a22o_2 _14326_ (.A1(\cpuregs[6][14] ),
    .A2(_11283_),
    .B1(_11290_),
    .B2(_11285_),
    .X(_03710_));
 sky130_fd_sc_hd__buf_1 _14327_ (.A(_11264_),
    .X(_11291_));
 sky130_fd_sc_hd__buf_1 _14328_ (.A(\cpuregs_wrdata[13] ),
    .X(_11292_));
 sky130_fd_sc_hd__buf_1 _14329_ (.A(_11268_),
    .X(_11293_));
 sky130_fd_sc_hd__a22o_2 _14330_ (.A1(\cpuregs[6][13] ),
    .A2(_11291_),
    .B1(_11292_),
    .B2(_11293_),
    .X(_03709_));
 sky130_fd_sc_hd__buf_1 _14331_ (.A(\cpuregs_wrdata[12] ),
    .X(_11294_));
 sky130_fd_sc_hd__a22o_2 _14332_ (.A1(\cpuregs[6][12] ),
    .A2(_11291_),
    .B1(_11294_),
    .B2(_11293_),
    .X(_03708_));
 sky130_fd_sc_hd__buf_1 _14333_ (.A(\cpuregs_wrdata[11] ),
    .X(_11295_));
 sky130_fd_sc_hd__a22o_2 _14334_ (.A1(\cpuregs[6][11] ),
    .A2(_11291_),
    .B1(_11295_),
    .B2(_11293_),
    .X(_03707_));
 sky130_fd_sc_hd__buf_1 _14335_ (.A(\cpuregs_wrdata[10] ),
    .X(_11296_));
 sky130_fd_sc_hd__a22o_2 _14336_ (.A1(\cpuregs[6][10] ),
    .A2(_11291_),
    .B1(_11296_),
    .B2(_11293_),
    .X(_03706_));
 sky130_fd_sc_hd__buf_1 _14337_ (.A(\cpuregs_wrdata[9] ),
    .X(_11297_));
 sky130_fd_sc_hd__a22o_2 _14338_ (.A1(\cpuregs[6][9] ),
    .A2(_11291_),
    .B1(_11297_),
    .B2(_11293_),
    .X(_03705_));
 sky130_fd_sc_hd__buf_1 _14339_ (.A(\cpuregs_wrdata[8] ),
    .X(_11298_));
 sky130_fd_sc_hd__a22o_2 _14340_ (.A1(\cpuregs[6][8] ),
    .A2(_11291_),
    .B1(_11298_),
    .B2(_11293_),
    .X(_03704_));
 sky130_fd_sc_hd__buf_1 _14341_ (.A(_11263_),
    .X(_11299_));
 sky130_fd_sc_hd__buf_1 _14342_ (.A(\cpuregs_wrdata[7] ),
    .X(_11300_));
 sky130_fd_sc_hd__buf_1 _14343_ (.A(_11267_),
    .X(_11301_));
 sky130_fd_sc_hd__a22o_2 _14344_ (.A1(\cpuregs[6][7] ),
    .A2(_11299_),
    .B1(_11300_),
    .B2(_11301_),
    .X(_03703_));
 sky130_fd_sc_hd__buf_1 _14345_ (.A(\cpuregs_wrdata[6] ),
    .X(_11302_));
 sky130_fd_sc_hd__a22o_2 _14346_ (.A1(\cpuregs[6][6] ),
    .A2(_11299_),
    .B1(_11302_),
    .B2(_11301_),
    .X(_03702_));
 sky130_fd_sc_hd__buf_1 _14347_ (.A(\cpuregs_wrdata[5] ),
    .X(_11303_));
 sky130_fd_sc_hd__a22o_2 _14348_ (.A1(\cpuregs[6][5] ),
    .A2(_11299_),
    .B1(_11303_),
    .B2(_11301_),
    .X(_03701_));
 sky130_fd_sc_hd__buf_1 _14349_ (.A(\cpuregs_wrdata[4] ),
    .X(_11304_));
 sky130_fd_sc_hd__a22o_2 _14350_ (.A1(\cpuregs[6][4] ),
    .A2(_11299_),
    .B1(_11304_),
    .B2(_11301_),
    .X(_03700_));
 sky130_fd_sc_hd__buf_1 _14351_ (.A(\cpuregs_wrdata[3] ),
    .X(_11305_));
 sky130_fd_sc_hd__a22o_2 _14352_ (.A1(\cpuregs[6][3] ),
    .A2(_11299_),
    .B1(_11305_),
    .B2(_11301_),
    .X(_03699_));
 sky130_fd_sc_hd__buf_1 _14353_ (.A(\cpuregs_wrdata[2] ),
    .X(_11306_));
 sky130_fd_sc_hd__a22o_2 _14354_ (.A1(\cpuregs[6][2] ),
    .A2(_11299_),
    .B1(_11306_),
    .B2(_11301_),
    .X(_03698_));
 sky130_fd_sc_hd__buf_1 _14355_ (.A(\cpuregs_wrdata[1] ),
    .X(_11307_));
 sky130_fd_sc_hd__a22o_2 _14356_ (.A1(\cpuregs[6][1] ),
    .A2(_11264_),
    .B1(_11307_),
    .B2(_11268_),
    .X(_03697_));
 sky130_fd_sc_hd__buf_1 _14357_ (.A(\cpuregs_wrdata[0] ),
    .X(_11308_));
 sky130_fd_sc_hd__a22o_2 _14358_ (.A1(\cpuregs[6][0] ),
    .A2(_11264_),
    .B1(_11308_),
    .B2(_11268_),
    .X(_03696_));
 sky130_vsdinv _14359_ (.A(\latched_rd[3] ),
    .Y(_11309_));
 sky130_fd_sc_hd__buf_1 _14360_ (.A(\latched_rd[2] ),
    .X(_11310_));
 sky130_fd_sc_hd__or3_2 _14361_ (.A(\latched_rd[4] ),
    .B(_11309_),
    .C(_11310_),
    .X(_11311_));
 sky130_vsdinv _14362_ (.A(\latched_rd[0] ),
    .Y(_11312_));
 sky130_fd_sc_hd__or3_2 _14363_ (.A(_11312_),
    .B(\latched_rd[1] ),
    .C(_11260_),
    .X(_11313_));
 sky130_fd_sc_hd__or2_2 _14364_ (.A(_11311_),
    .B(_11313_),
    .X(_11314_));
 sky130_fd_sc_hd__buf_1 _14365_ (.A(_11314_),
    .X(_11315_));
 sky130_fd_sc_hd__buf_1 _14366_ (.A(_11315_),
    .X(_11316_));
 sky130_vsdinv _14367_ (.A(_11314_),
    .Y(_11317_));
 sky130_fd_sc_hd__buf_1 _14368_ (.A(_11317_),
    .X(_11318_));
 sky130_fd_sc_hd__buf_1 _14369_ (.A(_11318_),
    .X(_11319_));
 sky130_fd_sc_hd__a22o_2 _14370_ (.A1(\cpuregs[9][31] ),
    .A2(_11316_),
    .B1(_11266_),
    .B2(_11319_),
    .X(_03695_));
 sky130_fd_sc_hd__a22o_2 _14371_ (.A1(\cpuregs[9][30] ),
    .A2(_11316_),
    .B1(_11270_),
    .B2(_11319_),
    .X(_03694_));
 sky130_fd_sc_hd__a22o_2 _14372_ (.A1(\cpuregs[9][29] ),
    .A2(_11316_),
    .B1(_11271_),
    .B2(_11319_),
    .X(_03693_));
 sky130_fd_sc_hd__a22o_2 _14373_ (.A1(\cpuregs[9][28] ),
    .A2(_11316_),
    .B1(_11272_),
    .B2(_11319_),
    .X(_03692_));
 sky130_fd_sc_hd__a22o_2 _14374_ (.A1(\cpuregs[9][27] ),
    .A2(_11316_),
    .B1(_11273_),
    .B2(_11319_),
    .X(_03691_));
 sky130_fd_sc_hd__a22o_2 _14375_ (.A1(\cpuregs[9][26] ),
    .A2(_11316_),
    .B1(_11274_),
    .B2(_11319_),
    .X(_03690_));
 sky130_fd_sc_hd__buf_1 _14376_ (.A(_11315_),
    .X(_11320_));
 sky130_fd_sc_hd__buf_1 _14377_ (.A(_11318_),
    .X(_11321_));
 sky130_fd_sc_hd__a22o_2 _14378_ (.A1(\cpuregs[9][25] ),
    .A2(_11320_),
    .B1(_11276_),
    .B2(_11321_),
    .X(_03689_));
 sky130_fd_sc_hd__a22o_2 _14379_ (.A1(\cpuregs[9][24] ),
    .A2(_11320_),
    .B1(_11278_),
    .B2(_11321_),
    .X(_03688_));
 sky130_fd_sc_hd__a22o_2 _14380_ (.A1(\cpuregs[9][23] ),
    .A2(_11320_),
    .B1(_11279_),
    .B2(_11321_),
    .X(_03687_));
 sky130_fd_sc_hd__a22o_2 _14381_ (.A1(\cpuregs[9][22] ),
    .A2(_11320_),
    .B1(_11280_),
    .B2(_11321_),
    .X(_03686_));
 sky130_fd_sc_hd__a22o_2 _14382_ (.A1(\cpuregs[9][21] ),
    .A2(_11320_),
    .B1(_11281_),
    .B2(_11321_),
    .X(_03685_));
 sky130_fd_sc_hd__a22o_2 _14383_ (.A1(\cpuregs[9][20] ),
    .A2(_11320_),
    .B1(_11282_),
    .B2(_11321_),
    .X(_03684_));
 sky130_fd_sc_hd__buf_1 _14384_ (.A(_11315_),
    .X(_11322_));
 sky130_fd_sc_hd__buf_1 _14385_ (.A(_11318_),
    .X(_11323_));
 sky130_fd_sc_hd__a22o_2 _14386_ (.A1(\cpuregs[9][19] ),
    .A2(_11322_),
    .B1(_11284_),
    .B2(_11323_),
    .X(_03683_));
 sky130_fd_sc_hd__a22o_2 _14387_ (.A1(\cpuregs[9][18] ),
    .A2(_11322_),
    .B1(_11286_),
    .B2(_11323_),
    .X(_03682_));
 sky130_fd_sc_hd__a22o_2 _14388_ (.A1(\cpuregs[9][17] ),
    .A2(_11322_),
    .B1(_11287_),
    .B2(_11323_),
    .X(_03681_));
 sky130_fd_sc_hd__a22o_2 _14389_ (.A1(\cpuregs[9][16] ),
    .A2(_11322_),
    .B1(_11288_),
    .B2(_11323_),
    .X(_03680_));
 sky130_fd_sc_hd__a22o_2 _14390_ (.A1(\cpuregs[9][15] ),
    .A2(_11322_),
    .B1(_11289_),
    .B2(_11323_),
    .X(_03679_));
 sky130_fd_sc_hd__a22o_2 _14391_ (.A1(\cpuregs[9][14] ),
    .A2(_11322_),
    .B1(_11290_),
    .B2(_11323_),
    .X(_03678_));
 sky130_fd_sc_hd__buf_1 _14392_ (.A(_11315_),
    .X(_11324_));
 sky130_fd_sc_hd__buf_1 _14393_ (.A(_11318_),
    .X(_11325_));
 sky130_fd_sc_hd__a22o_2 _14394_ (.A1(\cpuregs[9][13] ),
    .A2(_11324_),
    .B1(_11292_),
    .B2(_11325_),
    .X(_03677_));
 sky130_fd_sc_hd__a22o_2 _14395_ (.A1(\cpuregs[9][12] ),
    .A2(_11324_),
    .B1(_11294_),
    .B2(_11325_),
    .X(_03676_));
 sky130_fd_sc_hd__a22o_2 _14396_ (.A1(\cpuregs[9][11] ),
    .A2(_11324_),
    .B1(_11295_),
    .B2(_11325_),
    .X(_03675_));
 sky130_fd_sc_hd__a22o_2 _14397_ (.A1(\cpuregs[9][10] ),
    .A2(_11324_),
    .B1(_11296_),
    .B2(_11325_),
    .X(_03674_));
 sky130_fd_sc_hd__a22o_2 _14398_ (.A1(\cpuregs[9][9] ),
    .A2(_11324_),
    .B1(_11297_),
    .B2(_11325_),
    .X(_03673_));
 sky130_fd_sc_hd__a22o_2 _14399_ (.A1(\cpuregs[9][8] ),
    .A2(_11324_),
    .B1(_11298_),
    .B2(_11325_),
    .X(_03672_));
 sky130_fd_sc_hd__buf_1 _14400_ (.A(_11314_),
    .X(_11326_));
 sky130_fd_sc_hd__buf_1 _14401_ (.A(_11317_),
    .X(_11327_));
 sky130_fd_sc_hd__a22o_2 _14402_ (.A1(\cpuregs[9][7] ),
    .A2(_11326_),
    .B1(_11300_),
    .B2(_11327_),
    .X(_03671_));
 sky130_fd_sc_hd__a22o_2 _14403_ (.A1(\cpuregs[9][6] ),
    .A2(_11326_),
    .B1(_11302_),
    .B2(_11327_),
    .X(_03670_));
 sky130_fd_sc_hd__a22o_2 _14404_ (.A1(\cpuregs[9][5] ),
    .A2(_11326_),
    .B1(_11303_),
    .B2(_11327_),
    .X(_03669_));
 sky130_fd_sc_hd__a22o_2 _14405_ (.A1(\cpuregs[9][4] ),
    .A2(_11326_),
    .B1(_11304_),
    .B2(_11327_),
    .X(_03668_));
 sky130_fd_sc_hd__a22o_2 _14406_ (.A1(\cpuregs[9][3] ),
    .A2(_11326_),
    .B1(_11305_),
    .B2(_11327_),
    .X(_03667_));
 sky130_fd_sc_hd__a22o_2 _14407_ (.A1(\cpuregs[9][2] ),
    .A2(_11326_),
    .B1(_11306_),
    .B2(_11327_),
    .X(_03666_));
 sky130_fd_sc_hd__a22o_2 _14408_ (.A1(\cpuregs[9][1] ),
    .A2(_11315_),
    .B1(_11307_),
    .B2(_11318_),
    .X(_03665_));
 sky130_fd_sc_hd__a22o_2 _14409_ (.A1(\cpuregs[9][0] ),
    .A2(_11315_),
    .B1(_11308_),
    .B2(_11318_),
    .X(_03664_));
 sky130_fd_sc_hd__o21ai_2 _14410_ (.A1(\cpu_state[2] ),
    .A2(_10639_),
    .B1(_10443_),
    .Y(_11328_));
 sky130_fd_sc_hd__buf_1 _14411_ (.A(_11328_),
    .X(_11329_));
 sky130_fd_sc_hd__buf_1 _14412_ (.A(_11329_),
    .X(_11330_));
 sky130_vsdinv _14413_ (.A(_11328_),
    .Y(_11331_));
 sky130_fd_sc_hd__buf_1 _14414_ (.A(_11331_),
    .X(_11332_));
 sky130_fd_sc_hd__buf_1 _14415_ (.A(_11332_),
    .X(_11333_));
 sky130_fd_sc_hd__a22o_2 _14416_ (.A1(pcpi_rs2[31]),
    .A2(_11330_),
    .B1(_02467_),
    .B2(_11333_),
    .X(_03663_));
 sky130_fd_sc_hd__a22o_2 _14417_ (.A1(pcpi_rs2[30]),
    .A2(_11330_),
    .B1(_02466_),
    .B2(_11333_),
    .X(_03662_));
 sky130_fd_sc_hd__buf_1 _14418_ (.A(pcpi_rs2[29]),
    .X(_11334_));
 sky130_fd_sc_hd__a22o_2 _14419_ (.A1(_11334_),
    .A2(_11330_),
    .B1(_02464_),
    .B2(_11333_),
    .X(_03661_));
 sky130_fd_sc_hd__a22o_2 _14420_ (.A1(pcpi_rs2[28]),
    .A2(_11330_),
    .B1(_02463_),
    .B2(_11333_),
    .X(_03660_));
 sky130_fd_sc_hd__buf_1 _14421_ (.A(pcpi_rs2[27]),
    .X(_11335_));
 sky130_fd_sc_hd__a22o_2 _14422_ (.A1(_11335_),
    .A2(_11330_),
    .B1(_02462_),
    .B2(_11333_),
    .X(_03659_));
 sky130_fd_sc_hd__buf_1 _14423_ (.A(_11329_),
    .X(_11336_));
 sky130_fd_sc_hd__a22o_2 _14424_ (.A1(pcpi_rs2[26]),
    .A2(_11336_),
    .B1(_02461_),
    .B2(_11333_),
    .X(_03658_));
 sky130_fd_sc_hd__buf_1 _14425_ (.A(pcpi_rs2[25]),
    .X(_11337_));
 sky130_fd_sc_hd__buf_1 _14426_ (.A(_11332_),
    .X(_11338_));
 sky130_fd_sc_hd__a22o_2 _14427_ (.A1(_11337_),
    .A2(_11336_),
    .B1(_02460_),
    .B2(_11338_),
    .X(_03657_));
 sky130_fd_sc_hd__a22o_2 _14428_ (.A1(pcpi_rs2[24]),
    .A2(_11336_),
    .B1(_02459_),
    .B2(_11338_),
    .X(_03656_));
 sky130_fd_sc_hd__buf_1 _14429_ (.A(pcpi_rs2[23]),
    .X(_11339_));
 sky130_fd_sc_hd__a22o_2 _14430_ (.A1(_11339_),
    .A2(_11336_),
    .B1(_02458_),
    .B2(_11338_),
    .X(_03655_));
 sky130_fd_sc_hd__a22o_2 _14431_ (.A1(pcpi_rs2[22]),
    .A2(_11336_),
    .B1(_02457_),
    .B2(_11338_),
    .X(_03654_));
 sky130_fd_sc_hd__buf_1 _14432_ (.A(pcpi_rs2[21]),
    .X(_11340_));
 sky130_fd_sc_hd__a22o_2 _14433_ (.A1(_11340_),
    .A2(_11336_),
    .B1(_02456_),
    .B2(_11338_),
    .X(_03653_));
 sky130_fd_sc_hd__buf_1 _14434_ (.A(_11329_),
    .X(_11341_));
 sky130_fd_sc_hd__a22o_2 _14435_ (.A1(pcpi_rs2[20]),
    .A2(_11341_),
    .B1(_02455_),
    .B2(_11338_),
    .X(_03652_));
 sky130_fd_sc_hd__buf_1 _14436_ (.A(pcpi_rs2[19]),
    .X(_11342_));
 sky130_fd_sc_hd__buf_1 _14437_ (.A(_11332_),
    .X(_11343_));
 sky130_fd_sc_hd__a22o_2 _14438_ (.A1(_11342_),
    .A2(_11341_),
    .B1(_02453_),
    .B2(_11343_),
    .X(_03651_));
 sky130_fd_sc_hd__a22o_2 _14439_ (.A1(pcpi_rs2[18]),
    .A2(_11341_),
    .B1(_02452_),
    .B2(_11343_),
    .X(_03650_));
 sky130_fd_sc_hd__buf_1 _14440_ (.A(pcpi_rs2[17]),
    .X(_11344_));
 sky130_fd_sc_hd__a22o_2 _14441_ (.A1(_11344_),
    .A2(_11341_),
    .B1(_02451_),
    .B2(_11343_),
    .X(_03649_));
 sky130_fd_sc_hd__a22o_2 _14442_ (.A1(pcpi_rs2[16]),
    .A2(_11341_),
    .B1(_02450_),
    .B2(_11343_),
    .X(_03648_));
 sky130_fd_sc_hd__buf_1 _14443_ (.A(pcpi_rs2[15]),
    .X(_11345_));
 sky130_fd_sc_hd__a22o_2 _14444_ (.A1(_11345_),
    .A2(_11341_),
    .B1(_02449_),
    .B2(_11343_),
    .X(_03647_));
 sky130_fd_sc_hd__buf_1 _14445_ (.A(pcpi_rs2[14]),
    .X(_11346_));
 sky130_fd_sc_hd__buf_1 _14446_ (.A(_11328_),
    .X(_11347_));
 sky130_fd_sc_hd__a22o_2 _14447_ (.A1(_11346_),
    .A2(_11347_),
    .B1(_02448_),
    .B2(_11343_),
    .X(_03646_));
 sky130_fd_sc_hd__buf_1 _14448_ (.A(pcpi_rs2[13]),
    .X(_11348_));
 sky130_fd_sc_hd__buf_1 _14449_ (.A(_11332_),
    .X(_11349_));
 sky130_fd_sc_hd__a22o_2 _14450_ (.A1(_11348_),
    .A2(_11347_),
    .B1(_02447_),
    .B2(_11349_),
    .X(_03645_));
 sky130_fd_sc_hd__buf_1 _14451_ (.A(pcpi_rs2[12]),
    .X(_11350_));
 sky130_fd_sc_hd__a22o_2 _14452_ (.A1(_11350_),
    .A2(_11347_),
    .B1(_02446_),
    .B2(_11349_),
    .X(_03644_));
 sky130_fd_sc_hd__buf_1 _14453_ (.A(pcpi_rs2[11]),
    .X(_11351_));
 sky130_fd_sc_hd__a22o_2 _14454_ (.A1(_11351_),
    .A2(_11347_),
    .B1(_02445_),
    .B2(_11349_),
    .X(_03643_));
 sky130_fd_sc_hd__buf_1 _14455_ (.A(pcpi_rs2[10]),
    .X(_11352_));
 sky130_fd_sc_hd__a22o_2 _14456_ (.A1(_11352_),
    .A2(_11347_),
    .B1(_02444_),
    .B2(_11349_),
    .X(_03642_));
 sky130_fd_sc_hd__buf_1 _14457_ (.A(pcpi_rs2[9]),
    .X(_11353_));
 sky130_fd_sc_hd__a22o_2 _14458_ (.A1(_11353_),
    .A2(_11347_),
    .B1(_02474_),
    .B2(_11349_),
    .X(_03641_));
 sky130_fd_sc_hd__buf_1 _14459_ (.A(pcpi_rs2[8]),
    .X(_11354_));
 sky130_fd_sc_hd__buf_1 _14460_ (.A(_11328_),
    .X(_11355_));
 sky130_fd_sc_hd__a22o_2 _14461_ (.A1(_11354_),
    .A2(_11355_),
    .B1(_02473_),
    .B2(_11349_),
    .X(_03640_));
 sky130_fd_sc_hd__buf_1 _14462_ (.A(mem_la_wdata[7]),
    .X(_11356_));
 sky130_fd_sc_hd__buf_1 _14463_ (.A(_11331_),
    .X(_11357_));
 sky130_fd_sc_hd__a22o_2 _14464_ (.A1(_11356_),
    .A2(_11355_),
    .B1(_02472_),
    .B2(_11357_),
    .X(_03639_));
 sky130_fd_sc_hd__buf_1 _14465_ (.A(mem_la_wdata[6]),
    .X(_11358_));
 sky130_fd_sc_hd__a22o_2 _14466_ (.A1(_11358_),
    .A2(_11355_),
    .B1(_02471_),
    .B2(_11357_),
    .X(_03638_));
 sky130_fd_sc_hd__buf_1 _14467_ (.A(mem_la_wdata[5]),
    .X(_11359_));
 sky130_fd_sc_hd__a22o_2 _14468_ (.A1(_11359_),
    .A2(_11355_),
    .B1(_02470_),
    .B2(_11357_),
    .X(_03637_));
 sky130_fd_sc_hd__buf_1 _14469_ (.A(mem_la_wdata[4]),
    .X(_11360_));
 sky130_fd_sc_hd__a22o_2 _14470_ (.A1(_11360_),
    .A2(_11355_),
    .B1(_02469_),
    .B2(_11357_),
    .X(_03636_));
 sky130_fd_sc_hd__buf_1 _14471_ (.A(mem_la_wdata[3]),
    .X(_11361_));
 sky130_fd_sc_hd__a22o_2 _14472_ (.A1(_11361_),
    .A2(_11355_),
    .B1(_02468_),
    .B2(_11357_),
    .X(_03635_));
 sky130_fd_sc_hd__buf_1 _14473_ (.A(mem_la_wdata[2]),
    .X(_11362_));
 sky130_fd_sc_hd__a22o_2 _14474_ (.A1(_11362_),
    .A2(_11329_),
    .B1(_02465_),
    .B2(_11357_),
    .X(_03634_));
 sky130_fd_sc_hd__buf_1 _14475_ (.A(mem_la_wdata[1]),
    .X(_11363_));
 sky130_fd_sc_hd__a22o_2 _14476_ (.A1(_11363_),
    .A2(_11329_),
    .B1(_02454_),
    .B2(_11332_),
    .X(_03633_));
 sky130_fd_sc_hd__buf_1 _14477_ (.A(mem_la_wdata[0]),
    .X(_11364_));
 sky130_fd_sc_hd__a22o_2 _14478_ (.A1(_11364_),
    .A2(_11329_),
    .B1(_02443_),
    .B2(_11332_),
    .X(_03632_));
 sky130_fd_sc_hd__or3_2 _14479_ (.A(\latched_rd[0] ),
    .B(\latched_rd[1] ),
    .C(_11260_),
    .X(_11365_));
 sky130_fd_sc_hd__or2_2 _14480_ (.A(_11254_),
    .B(_11365_),
    .X(_11366_));
 sky130_fd_sc_hd__buf_1 _14481_ (.A(_11366_),
    .X(_11367_));
 sky130_fd_sc_hd__buf_1 _14482_ (.A(_11367_),
    .X(_11368_));
 sky130_vsdinv _14483_ (.A(_11366_),
    .Y(_11369_));
 sky130_fd_sc_hd__buf_1 _14484_ (.A(_11369_),
    .X(_11370_));
 sky130_fd_sc_hd__buf_1 _14485_ (.A(_11370_),
    .X(_11371_));
 sky130_fd_sc_hd__a22o_2 _14486_ (.A1(\cpuregs[4][31] ),
    .A2(_11368_),
    .B1(_11266_),
    .B2(_11371_),
    .X(_03631_));
 sky130_fd_sc_hd__a22o_2 _14487_ (.A1(\cpuregs[4][30] ),
    .A2(_11368_),
    .B1(_11270_),
    .B2(_11371_),
    .X(_03630_));
 sky130_fd_sc_hd__a22o_2 _14488_ (.A1(\cpuregs[4][29] ),
    .A2(_11368_),
    .B1(_11271_),
    .B2(_11371_),
    .X(_03629_));
 sky130_fd_sc_hd__a22o_2 _14489_ (.A1(\cpuregs[4][28] ),
    .A2(_11368_),
    .B1(_11272_),
    .B2(_11371_),
    .X(_03628_));
 sky130_fd_sc_hd__a22o_2 _14490_ (.A1(\cpuregs[4][27] ),
    .A2(_11368_),
    .B1(_11273_),
    .B2(_11371_),
    .X(_03627_));
 sky130_fd_sc_hd__a22o_2 _14491_ (.A1(\cpuregs[4][26] ),
    .A2(_11368_),
    .B1(_11274_),
    .B2(_11371_),
    .X(_03626_));
 sky130_fd_sc_hd__buf_1 _14492_ (.A(_11367_),
    .X(_11372_));
 sky130_fd_sc_hd__buf_1 _14493_ (.A(_11370_),
    .X(_11373_));
 sky130_fd_sc_hd__a22o_2 _14494_ (.A1(\cpuregs[4][25] ),
    .A2(_11372_),
    .B1(_11276_),
    .B2(_11373_),
    .X(_03625_));
 sky130_fd_sc_hd__a22o_2 _14495_ (.A1(\cpuregs[4][24] ),
    .A2(_11372_),
    .B1(_11278_),
    .B2(_11373_),
    .X(_03624_));
 sky130_fd_sc_hd__a22o_2 _14496_ (.A1(\cpuregs[4][23] ),
    .A2(_11372_),
    .B1(_11279_),
    .B2(_11373_),
    .X(_03623_));
 sky130_fd_sc_hd__a22o_2 _14497_ (.A1(\cpuregs[4][22] ),
    .A2(_11372_),
    .B1(_11280_),
    .B2(_11373_),
    .X(_03622_));
 sky130_fd_sc_hd__a22o_2 _14498_ (.A1(\cpuregs[4][21] ),
    .A2(_11372_),
    .B1(_11281_),
    .B2(_11373_),
    .X(_03621_));
 sky130_fd_sc_hd__a22o_2 _14499_ (.A1(\cpuregs[4][20] ),
    .A2(_11372_),
    .B1(_11282_),
    .B2(_11373_),
    .X(_03620_));
 sky130_fd_sc_hd__buf_1 _14500_ (.A(_11367_),
    .X(_11374_));
 sky130_fd_sc_hd__buf_1 _14501_ (.A(_11370_),
    .X(_11375_));
 sky130_fd_sc_hd__a22o_2 _14502_ (.A1(\cpuregs[4][19] ),
    .A2(_11374_),
    .B1(_11284_),
    .B2(_11375_),
    .X(_03619_));
 sky130_fd_sc_hd__a22o_2 _14503_ (.A1(\cpuregs[4][18] ),
    .A2(_11374_),
    .B1(_11286_),
    .B2(_11375_),
    .X(_03618_));
 sky130_fd_sc_hd__a22o_2 _14504_ (.A1(\cpuregs[4][17] ),
    .A2(_11374_),
    .B1(_11287_),
    .B2(_11375_),
    .X(_03617_));
 sky130_fd_sc_hd__a22o_2 _14505_ (.A1(\cpuregs[4][16] ),
    .A2(_11374_),
    .B1(_11288_),
    .B2(_11375_),
    .X(_03616_));
 sky130_fd_sc_hd__a22o_2 _14506_ (.A1(\cpuregs[4][15] ),
    .A2(_11374_),
    .B1(_11289_),
    .B2(_11375_),
    .X(_03615_));
 sky130_fd_sc_hd__a22o_2 _14507_ (.A1(\cpuregs[4][14] ),
    .A2(_11374_),
    .B1(_11290_),
    .B2(_11375_),
    .X(_03614_));
 sky130_fd_sc_hd__buf_1 _14508_ (.A(_11367_),
    .X(_11376_));
 sky130_fd_sc_hd__buf_1 _14509_ (.A(_11370_),
    .X(_11377_));
 sky130_fd_sc_hd__a22o_2 _14510_ (.A1(\cpuregs[4][13] ),
    .A2(_11376_),
    .B1(_11292_),
    .B2(_11377_),
    .X(_03613_));
 sky130_fd_sc_hd__a22o_2 _14511_ (.A1(\cpuregs[4][12] ),
    .A2(_11376_),
    .B1(_11294_),
    .B2(_11377_),
    .X(_03612_));
 sky130_fd_sc_hd__a22o_2 _14512_ (.A1(\cpuregs[4][11] ),
    .A2(_11376_),
    .B1(_11295_),
    .B2(_11377_),
    .X(_03611_));
 sky130_fd_sc_hd__a22o_2 _14513_ (.A1(\cpuregs[4][10] ),
    .A2(_11376_),
    .B1(_11296_),
    .B2(_11377_),
    .X(_03610_));
 sky130_fd_sc_hd__a22o_2 _14514_ (.A1(\cpuregs[4][9] ),
    .A2(_11376_),
    .B1(_11297_),
    .B2(_11377_),
    .X(_03609_));
 sky130_fd_sc_hd__a22o_2 _14515_ (.A1(\cpuregs[4][8] ),
    .A2(_11376_),
    .B1(_11298_),
    .B2(_11377_),
    .X(_03608_));
 sky130_fd_sc_hd__buf_1 _14516_ (.A(_11366_),
    .X(_11378_));
 sky130_fd_sc_hd__buf_1 _14517_ (.A(_11369_),
    .X(_11379_));
 sky130_fd_sc_hd__a22o_2 _14518_ (.A1(\cpuregs[4][7] ),
    .A2(_11378_),
    .B1(_11300_),
    .B2(_11379_),
    .X(_03607_));
 sky130_fd_sc_hd__a22o_2 _14519_ (.A1(\cpuregs[4][6] ),
    .A2(_11378_),
    .B1(_11302_),
    .B2(_11379_),
    .X(_03606_));
 sky130_fd_sc_hd__a22o_2 _14520_ (.A1(\cpuregs[4][5] ),
    .A2(_11378_),
    .B1(_11303_),
    .B2(_11379_),
    .X(_03605_));
 sky130_fd_sc_hd__a22o_2 _14521_ (.A1(\cpuregs[4][4] ),
    .A2(_11378_),
    .B1(_11304_),
    .B2(_11379_),
    .X(_03604_));
 sky130_fd_sc_hd__a22o_2 _14522_ (.A1(\cpuregs[4][3] ),
    .A2(_11378_),
    .B1(_11305_),
    .B2(_11379_),
    .X(_03603_));
 sky130_fd_sc_hd__a22o_2 _14523_ (.A1(\cpuregs[4][2] ),
    .A2(_11378_),
    .B1(_11306_),
    .B2(_11379_),
    .X(_03602_));
 sky130_fd_sc_hd__a22o_2 _14524_ (.A1(\cpuregs[4][1] ),
    .A2(_11367_),
    .B1(_11307_),
    .B2(_11370_),
    .X(_03601_));
 sky130_fd_sc_hd__a22o_2 _14525_ (.A1(\cpuregs[4][0] ),
    .A2(_11367_),
    .B1(_11308_),
    .B2(_11370_),
    .X(_03600_));
 sky130_vsdinv _14526_ (.A(\latched_rd[4] ),
    .Y(_11380_));
 sky130_fd_sc_hd__or2_2 _14527_ (.A(_11312_),
    .B(_11261_),
    .X(_11381_));
 sky130_fd_sc_hd__or4_2 _14528_ (.A(_11380_),
    .B(_11310_),
    .C(_11252_),
    .D(_11381_),
    .X(_11382_));
 sky130_fd_sc_hd__buf_1 _14529_ (.A(_11382_),
    .X(_11383_));
 sky130_fd_sc_hd__buf_1 _14530_ (.A(_11383_),
    .X(_11384_));
 sky130_vsdinv _14531_ (.A(_11382_),
    .Y(_11385_));
 sky130_fd_sc_hd__buf_1 _14532_ (.A(_11385_),
    .X(_11386_));
 sky130_fd_sc_hd__buf_1 _14533_ (.A(_11386_),
    .X(_11387_));
 sky130_fd_sc_hd__a22o_2 _14534_ (.A1(\cpuregs[19][31] ),
    .A2(_11384_),
    .B1(_11266_),
    .B2(_11387_),
    .X(_03599_));
 sky130_fd_sc_hd__a22o_2 _14535_ (.A1(\cpuregs[19][30] ),
    .A2(_11384_),
    .B1(_11270_),
    .B2(_11387_),
    .X(_03598_));
 sky130_fd_sc_hd__a22o_2 _14536_ (.A1(\cpuregs[19][29] ),
    .A2(_11384_),
    .B1(_11271_),
    .B2(_11387_),
    .X(_03597_));
 sky130_fd_sc_hd__a22o_2 _14537_ (.A1(\cpuregs[19][28] ),
    .A2(_11384_),
    .B1(_11272_),
    .B2(_11387_),
    .X(_03596_));
 sky130_fd_sc_hd__a22o_2 _14538_ (.A1(\cpuregs[19][27] ),
    .A2(_11384_),
    .B1(_11273_),
    .B2(_11387_),
    .X(_03595_));
 sky130_fd_sc_hd__a22o_2 _14539_ (.A1(\cpuregs[19][26] ),
    .A2(_11384_),
    .B1(_11274_),
    .B2(_11387_),
    .X(_03594_));
 sky130_fd_sc_hd__buf_1 _14540_ (.A(_11383_),
    .X(_11388_));
 sky130_fd_sc_hd__buf_1 _14541_ (.A(_11386_),
    .X(_11389_));
 sky130_fd_sc_hd__a22o_2 _14542_ (.A1(\cpuregs[19][25] ),
    .A2(_11388_),
    .B1(_11276_),
    .B2(_11389_),
    .X(_03593_));
 sky130_fd_sc_hd__a22o_2 _14543_ (.A1(\cpuregs[19][24] ),
    .A2(_11388_),
    .B1(_11278_),
    .B2(_11389_),
    .X(_03592_));
 sky130_fd_sc_hd__a22o_2 _14544_ (.A1(\cpuregs[19][23] ),
    .A2(_11388_),
    .B1(_11279_),
    .B2(_11389_),
    .X(_03591_));
 sky130_fd_sc_hd__a22o_2 _14545_ (.A1(\cpuregs[19][22] ),
    .A2(_11388_),
    .B1(_11280_),
    .B2(_11389_),
    .X(_03590_));
 sky130_fd_sc_hd__a22o_2 _14546_ (.A1(\cpuregs[19][21] ),
    .A2(_11388_),
    .B1(_11281_),
    .B2(_11389_),
    .X(_03589_));
 sky130_fd_sc_hd__a22o_2 _14547_ (.A1(\cpuregs[19][20] ),
    .A2(_11388_),
    .B1(_11282_),
    .B2(_11389_),
    .X(_03588_));
 sky130_fd_sc_hd__buf_1 _14548_ (.A(_11383_),
    .X(_11390_));
 sky130_fd_sc_hd__buf_1 _14549_ (.A(_11386_),
    .X(_11391_));
 sky130_fd_sc_hd__a22o_2 _14550_ (.A1(\cpuregs[19][19] ),
    .A2(_11390_),
    .B1(_11284_),
    .B2(_11391_),
    .X(_03587_));
 sky130_fd_sc_hd__a22o_2 _14551_ (.A1(\cpuregs[19][18] ),
    .A2(_11390_),
    .B1(_11286_),
    .B2(_11391_),
    .X(_03586_));
 sky130_fd_sc_hd__a22o_2 _14552_ (.A1(\cpuregs[19][17] ),
    .A2(_11390_),
    .B1(_11287_),
    .B2(_11391_),
    .X(_03585_));
 sky130_fd_sc_hd__a22o_2 _14553_ (.A1(\cpuregs[19][16] ),
    .A2(_11390_),
    .B1(_11288_),
    .B2(_11391_),
    .X(_03584_));
 sky130_fd_sc_hd__a22o_2 _14554_ (.A1(\cpuregs[19][15] ),
    .A2(_11390_),
    .B1(_11289_),
    .B2(_11391_),
    .X(_03583_));
 sky130_fd_sc_hd__a22o_2 _14555_ (.A1(\cpuregs[19][14] ),
    .A2(_11390_),
    .B1(_11290_),
    .B2(_11391_),
    .X(_03582_));
 sky130_fd_sc_hd__buf_1 _14556_ (.A(_11383_),
    .X(_11392_));
 sky130_fd_sc_hd__buf_1 _14557_ (.A(_11386_),
    .X(_11393_));
 sky130_fd_sc_hd__a22o_2 _14558_ (.A1(\cpuregs[19][13] ),
    .A2(_11392_),
    .B1(_11292_),
    .B2(_11393_),
    .X(_03581_));
 sky130_fd_sc_hd__a22o_2 _14559_ (.A1(\cpuregs[19][12] ),
    .A2(_11392_),
    .B1(_11294_),
    .B2(_11393_),
    .X(_03580_));
 sky130_fd_sc_hd__a22o_2 _14560_ (.A1(\cpuregs[19][11] ),
    .A2(_11392_),
    .B1(_11295_),
    .B2(_11393_),
    .X(_03579_));
 sky130_fd_sc_hd__a22o_2 _14561_ (.A1(\cpuregs[19][10] ),
    .A2(_11392_),
    .B1(_11296_),
    .B2(_11393_),
    .X(_03578_));
 sky130_fd_sc_hd__a22o_2 _14562_ (.A1(\cpuregs[19][9] ),
    .A2(_11392_),
    .B1(_11297_),
    .B2(_11393_),
    .X(_03577_));
 sky130_fd_sc_hd__a22o_2 _14563_ (.A1(\cpuregs[19][8] ),
    .A2(_11392_),
    .B1(_11298_),
    .B2(_11393_),
    .X(_03576_));
 sky130_fd_sc_hd__buf_1 _14564_ (.A(_11382_),
    .X(_11394_));
 sky130_fd_sc_hd__buf_1 _14565_ (.A(_11385_),
    .X(_11395_));
 sky130_fd_sc_hd__a22o_2 _14566_ (.A1(\cpuregs[19][7] ),
    .A2(_11394_),
    .B1(_11300_),
    .B2(_11395_),
    .X(_03575_));
 sky130_fd_sc_hd__a22o_2 _14567_ (.A1(\cpuregs[19][6] ),
    .A2(_11394_),
    .B1(_11302_),
    .B2(_11395_),
    .X(_03574_));
 sky130_fd_sc_hd__a22o_2 _14568_ (.A1(\cpuregs[19][5] ),
    .A2(_11394_),
    .B1(_11303_),
    .B2(_11395_),
    .X(_03573_));
 sky130_fd_sc_hd__a22o_2 _14569_ (.A1(\cpuregs[19][4] ),
    .A2(_11394_),
    .B1(_11304_),
    .B2(_11395_),
    .X(_03572_));
 sky130_fd_sc_hd__a22o_2 _14570_ (.A1(\cpuregs[19][3] ),
    .A2(_11394_),
    .B1(_11305_),
    .B2(_11395_),
    .X(_03571_));
 sky130_fd_sc_hd__a22o_2 _14571_ (.A1(\cpuregs[19][2] ),
    .A2(_11394_),
    .B1(_11306_),
    .B2(_11395_),
    .X(_03570_));
 sky130_fd_sc_hd__a22o_2 _14572_ (.A1(\cpuregs[19][1] ),
    .A2(_11383_),
    .B1(_11307_),
    .B2(_11386_),
    .X(_03569_));
 sky130_fd_sc_hd__a22o_2 _14573_ (.A1(\cpuregs[19][0] ),
    .A2(_11383_),
    .B1(_11308_),
    .B2(_11386_),
    .X(_03568_));
 sky130_fd_sc_hd__or3_2 _14574_ (.A(_10475_),
    .B(_10452_),
    .C(_10708_),
    .X(_11396_));
 sky130_fd_sc_hd__or2_2 _14575_ (.A(trap),
    .B(_11396_),
    .X(_11397_));
 sky130_fd_sc_hd__buf_1 _14576_ (.A(_11397_),
    .X(_11398_));
 sky130_fd_sc_hd__buf_1 _14577_ (.A(_11398_),
    .X(_11399_));
 sky130_vsdinv _14578_ (.A(_11397_),
    .Y(_11400_));
 sky130_fd_sc_hd__buf_1 _14579_ (.A(_11400_),
    .X(_11401_));
 sky130_fd_sc_hd__buf_1 _14580_ (.A(_11401_),
    .X(_11402_));
 sky130_fd_sc_hd__a22o_2 _14581_ (.A1(mem_wdata[31]),
    .A2(_11399_),
    .B1(mem_la_wdata[31]),
    .B2(_11402_),
    .X(_03567_));
 sky130_fd_sc_hd__a22o_2 _14582_ (.A1(mem_wdata[30]),
    .A2(_11399_),
    .B1(mem_la_wdata[30]),
    .B2(_11402_),
    .X(_03566_));
 sky130_fd_sc_hd__a22o_2 _14583_ (.A1(mem_wdata[29]),
    .A2(_11399_),
    .B1(mem_la_wdata[29]),
    .B2(_11402_),
    .X(_03565_));
 sky130_fd_sc_hd__a22o_2 _14584_ (.A1(mem_wdata[28]),
    .A2(_11399_),
    .B1(mem_la_wdata[28]),
    .B2(_11402_),
    .X(_03564_));
 sky130_fd_sc_hd__a22o_2 _14585_ (.A1(mem_wdata[27]),
    .A2(_11399_),
    .B1(mem_la_wdata[27]),
    .B2(_11402_),
    .X(_03563_));
 sky130_fd_sc_hd__a22o_2 _14586_ (.A1(mem_wdata[26]),
    .A2(_11399_),
    .B1(mem_la_wdata[26]),
    .B2(_11402_),
    .X(_03562_));
 sky130_fd_sc_hd__buf_1 _14587_ (.A(_11398_),
    .X(_11403_));
 sky130_fd_sc_hd__buf_1 _14588_ (.A(_11401_),
    .X(_11404_));
 sky130_fd_sc_hd__a22o_2 _14589_ (.A1(mem_wdata[25]),
    .A2(_11403_),
    .B1(mem_la_wdata[25]),
    .B2(_11404_),
    .X(_03561_));
 sky130_fd_sc_hd__a22o_2 _14590_ (.A1(mem_wdata[24]),
    .A2(_11403_),
    .B1(mem_la_wdata[24]),
    .B2(_11404_),
    .X(_03560_));
 sky130_fd_sc_hd__a22o_2 _14591_ (.A1(mem_wdata[23]),
    .A2(_11403_),
    .B1(mem_la_wdata[23]),
    .B2(_11404_),
    .X(_03559_));
 sky130_fd_sc_hd__a22o_2 _14592_ (.A1(mem_wdata[22]),
    .A2(_11403_),
    .B1(mem_la_wdata[22]),
    .B2(_11404_),
    .X(_03558_));
 sky130_fd_sc_hd__a22o_2 _14593_ (.A1(mem_wdata[21]),
    .A2(_11403_),
    .B1(mem_la_wdata[21]),
    .B2(_11404_),
    .X(_03557_));
 sky130_fd_sc_hd__a22o_2 _14594_ (.A1(mem_wdata[20]),
    .A2(_11403_),
    .B1(mem_la_wdata[20]),
    .B2(_11404_),
    .X(_03556_));
 sky130_fd_sc_hd__buf_1 _14595_ (.A(_11398_),
    .X(_11405_));
 sky130_fd_sc_hd__buf_1 _14596_ (.A(_11401_),
    .X(_11406_));
 sky130_fd_sc_hd__a22o_2 _14597_ (.A1(mem_wdata[19]),
    .A2(_11405_),
    .B1(mem_la_wdata[19]),
    .B2(_11406_),
    .X(_03555_));
 sky130_fd_sc_hd__a22o_2 _14598_ (.A1(mem_wdata[18]),
    .A2(_11405_),
    .B1(mem_la_wdata[18]),
    .B2(_11406_),
    .X(_03554_));
 sky130_fd_sc_hd__a22o_2 _14599_ (.A1(mem_wdata[17]),
    .A2(_11405_),
    .B1(mem_la_wdata[17]),
    .B2(_11406_),
    .X(_03553_));
 sky130_fd_sc_hd__a22o_2 _14600_ (.A1(mem_wdata[16]),
    .A2(_11405_),
    .B1(mem_la_wdata[16]),
    .B2(_11406_),
    .X(_03552_));
 sky130_fd_sc_hd__a22o_2 _14601_ (.A1(mem_wdata[15]),
    .A2(_11405_),
    .B1(mem_la_wdata[15]),
    .B2(_11406_),
    .X(_03551_));
 sky130_fd_sc_hd__a22o_2 _14602_ (.A1(mem_wdata[14]),
    .A2(_11405_),
    .B1(mem_la_wdata[14]),
    .B2(_11406_),
    .X(_03550_));
 sky130_fd_sc_hd__buf_1 _14603_ (.A(_11398_),
    .X(_11407_));
 sky130_fd_sc_hd__buf_1 _14604_ (.A(_11401_),
    .X(_11408_));
 sky130_fd_sc_hd__a22o_2 _14605_ (.A1(mem_wdata[13]),
    .A2(_11407_),
    .B1(mem_la_wdata[13]),
    .B2(_11408_),
    .X(_03549_));
 sky130_fd_sc_hd__a22o_2 _14606_ (.A1(mem_wdata[12]),
    .A2(_11407_),
    .B1(mem_la_wdata[12]),
    .B2(_11408_),
    .X(_03548_));
 sky130_fd_sc_hd__a22o_2 _14607_ (.A1(mem_wdata[11]),
    .A2(_11407_),
    .B1(mem_la_wdata[11]),
    .B2(_11408_),
    .X(_03547_));
 sky130_fd_sc_hd__a22o_2 _14608_ (.A1(mem_wdata[10]),
    .A2(_11407_),
    .B1(mem_la_wdata[10]),
    .B2(_11408_),
    .X(_03546_));
 sky130_fd_sc_hd__a22o_2 _14609_ (.A1(mem_wdata[9]),
    .A2(_11407_),
    .B1(mem_la_wdata[9]),
    .B2(_11408_),
    .X(_03545_));
 sky130_fd_sc_hd__a22o_2 _14610_ (.A1(mem_wdata[8]),
    .A2(_11407_),
    .B1(mem_la_wdata[8]),
    .B2(_11408_),
    .X(_03544_));
 sky130_fd_sc_hd__buf_1 _14611_ (.A(_11397_),
    .X(_11409_));
 sky130_fd_sc_hd__buf_1 _14612_ (.A(_11400_),
    .X(_11410_));
 sky130_fd_sc_hd__a22o_2 _14613_ (.A1(mem_wdata[7]),
    .A2(_11409_),
    .B1(_11356_),
    .B2(_11410_),
    .X(_03543_));
 sky130_fd_sc_hd__a22o_2 _14614_ (.A1(mem_wdata[6]),
    .A2(_11409_),
    .B1(_11358_),
    .B2(_11410_),
    .X(_03542_));
 sky130_fd_sc_hd__a22o_2 _14615_ (.A1(mem_wdata[5]),
    .A2(_11409_),
    .B1(_11359_),
    .B2(_11410_),
    .X(_03541_));
 sky130_fd_sc_hd__a22o_2 _14616_ (.A1(mem_wdata[4]),
    .A2(_11409_),
    .B1(_11360_),
    .B2(_11410_),
    .X(_03540_));
 sky130_fd_sc_hd__a22o_2 _14617_ (.A1(mem_wdata[3]),
    .A2(_11409_),
    .B1(_11361_),
    .B2(_11410_),
    .X(_03539_));
 sky130_fd_sc_hd__a22o_2 _14618_ (.A1(mem_wdata[2]),
    .A2(_11409_),
    .B1(_11362_),
    .B2(_11410_),
    .X(_03538_));
 sky130_fd_sc_hd__a22o_2 _14619_ (.A1(mem_wdata[1]),
    .A2(_11398_),
    .B1(_11363_),
    .B2(_11401_),
    .X(_03537_));
 sky130_fd_sc_hd__a22o_2 _14620_ (.A1(mem_wdata[0]),
    .A2(_11398_),
    .B1(_11364_),
    .B2(_11401_),
    .X(_03536_));
 sky130_fd_sc_hd__or2_2 _14621_ (.A(_11254_),
    .B(_11381_),
    .X(_11411_));
 sky130_fd_sc_hd__buf_1 _14622_ (.A(_11411_),
    .X(_11412_));
 sky130_fd_sc_hd__buf_1 _14623_ (.A(_11412_),
    .X(_11413_));
 sky130_vsdinv _14624_ (.A(_11411_),
    .Y(_11414_));
 sky130_fd_sc_hd__buf_1 _14625_ (.A(_11414_),
    .X(_11415_));
 sky130_fd_sc_hd__buf_1 _14626_ (.A(_11415_),
    .X(_11416_));
 sky130_fd_sc_hd__a22o_2 _14627_ (.A1(\cpuregs[7][31] ),
    .A2(_11413_),
    .B1(_11266_),
    .B2(_11416_),
    .X(_03535_));
 sky130_fd_sc_hd__a22o_2 _14628_ (.A1(\cpuregs[7][30] ),
    .A2(_11413_),
    .B1(_11270_),
    .B2(_11416_),
    .X(_03534_));
 sky130_fd_sc_hd__a22o_2 _14629_ (.A1(\cpuregs[7][29] ),
    .A2(_11413_),
    .B1(_11271_),
    .B2(_11416_),
    .X(_03533_));
 sky130_fd_sc_hd__a22o_2 _14630_ (.A1(\cpuregs[7][28] ),
    .A2(_11413_),
    .B1(_11272_),
    .B2(_11416_),
    .X(_03532_));
 sky130_fd_sc_hd__a22o_2 _14631_ (.A1(\cpuregs[7][27] ),
    .A2(_11413_),
    .B1(_11273_),
    .B2(_11416_),
    .X(_03531_));
 sky130_fd_sc_hd__a22o_2 _14632_ (.A1(\cpuregs[7][26] ),
    .A2(_11413_),
    .B1(_11274_),
    .B2(_11416_),
    .X(_03530_));
 sky130_fd_sc_hd__buf_1 _14633_ (.A(_11412_),
    .X(_11417_));
 sky130_fd_sc_hd__buf_1 _14634_ (.A(_11415_),
    .X(_11418_));
 sky130_fd_sc_hd__a22o_2 _14635_ (.A1(\cpuregs[7][25] ),
    .A2(_11417_),
    .B1(_11276_),
    .B2(_11418_),
    .X(_03529_));
 sky130_fd_sc_hd__a22o_2 _14636_ (.A1(\cpuregs[7][24] ),
    .A2(_11417_),
    .B1(_11278_),
    .B2(_11418_),
    .X(_03528_));
 sky130_fd_sc_hd__a22o_2 _14637_ (.A1(\cpuregs[7][23] ),
    .A2(_11417_),
    .B1(_11279_),
    .B2(_11418_),
    .X(_03527_));
 sky130_fd_sc_hd__a22o_2 _14638_ (.A1(\cpuregs[7][22] ),
    .A2(_11417_),
    .B1(_11280_),
    .B2(_11418_),
    .X(_03526_));
 sky130_fd_sc_hd__a22o_2 _14639_ (.A1(\cpuregs[7][21] ),
    .A2(_11417_),
    .B1(_11281_),
    .B2(_11418_),
    .X(_03525_));
 sky130_fd_sc_hd__a22o_2 _14640_ (.A1(\cpuregs[7][20] ),
    .A2(_11417_),
    .B1(_11282_),
    .B2(_11418_),
    .X(_03524_));
 sky130_fd_sc_hd__buf_1 _14641_ (.A(_11412_),
    .X(_11419_));
 sky130_fd_sc_hd__buf_1 _14642_ (.A(_11415_),
    .X(_11420_));
 sky130_fd_sc_hd__a22o_2 _14643_ (.A1(\cpuregs[7][19] ),
    .A2(_11419_),
    .B1(_11284_),
    .B2(_11420_),
    .X(_03523_));
 sky130_fd_sc_hd__a22o_2 _14644_ (.A1(\cpuregs[7][18] ),
    .A2(_11419_),
    .B1(_11286_),
    .B2(_11420_),
    .X(_03522_));
 sky130_fd_sc_hd__a22o_2 _14645_ (.A1(\cpuregs[7][17] ),
    .A2(_11419_),
    .B1(_11287_),
    .B2(_11420_),
    .X(_03521_));
 sky130_fd_sc_hd__a22o_2 _14646_ (.A1(\cpuregs[7][16] ),
    .A2(_11419_),
    .B1(_11288_),
    .B2(_11420_),
    .X(_03520_));
 sky130_fd_sc_hd__a22o_2 _14647_ (.A1(\cpuregs[7][15] ),
    .A2(_11419_),
    .B1(_11289_),
    .B2(_11420_),
    .X(_03519_));
 sky130_fd_sc_hd__a22o_2 _14648_ (.A1(\cpuregs[7][14] ),
    .A2(_11419_),
    .B1(_11290_),
    .B2(_11420_),
    .X(_03518_));
 sky130_fd_sc_hd__buf_1 _14649_ (.A(_11412_),
    .X(_11421_));
 sky130_fd_sc_hd__buf_1 _14650_ (.A(_11415_),
    .X(_11422_));
 sky130_fd_sc_hd__a22o_2 _14651_ (.A1(\cpuregs[7][13] ),
    .A2(_11421_),
    .B1(_11292_),
    .B2(_11422_),
    .X(_03517_));
 sky130_fd_sc_hd__a22o_2 _14652_ (.A1(\cpuregs[7][12] ),
    .A2(_11421_),
    .B1(_11294_),
    .B2(_11422_),
    .X(_03516_));
 sky130_fd_sc_hd__a22o_2 _14653_ (.A1(\cpuregs[7][11] ),
    .A2(_11421_),
    .B1(_11295_),
    .B2(_11422_),
    .X(_03515_));
 sky130_fd_sc_hd__a22o_2 _14654_ (.A1(\cpuregs[7][10] ),
    .A2(_11421_),
    .B1(_11296_),
    .B2(_11422_),
    .X(_03514_));
 sky130_fd_sc_hd__a22o_2 _14655_ (.A1(\cpuregs[7][9] ),
    .A2(_11421_),
    .B1(_11297_),
    .B2(_11422_),
    .X(_03513_));
 sky130_fd_sc_hd__a22o_2 _14656_ (.A1(\cpuregs[7][8] ),
    .A2(_11421_),
    .B1(_11298_),
    .B2(_11422_),
    .X(_03512_));
 sky130_fd_sc_hd__buf_1 _14657_ (.A(_11411_),
    .X(_11423_));
 sky130_fd_sc_hd__buf_1 _14658_ (.A(_11414_),
    .X(_11424_));
 sky130_fd_sc_hd__a22o_2 _14659_ (.A1(\cpuregs[7][7] ),
    .A2(_11423_),
    .B1(_11300_),
    .B2(_11424_),
    .X(_03511_));
 sky130_fd_sc_hd__a22o_2 _14660_ (.A1(\cpuregs[7][6] ),
    .A2(_11423_),
    .B1(_11302_),
    .B2(_11424_),
    .X(_03510_));
 sky130_fd_sc_hd__a22o_2 _14661_ (.A1(\cpuregs[7][5] ),
    .A2(_11423_),
    .B1(_11303_),
    .B2(_11424_),
    .X(_03509_));
 sky130_fd_sc_hd__a22o_2 _14662_ (.A1(\cpuregs[7][4] ),
    .A2(_11423_),
    .B1(_11304_),
    .B2(_11424_),
    .X(_03508_));
 sky130_fd_sc_hd__a22o_2 _14663_ (.A1(\cpuregs[7][3] ),
    .A2(_11423_),
    .B1(_11305_),
    .B2(_11424_),
    .X(_03507_));
 sky130_fd_sc_hd__a22o_2 _14664_ (.A1(\cpuregs[7][2] ),
    .A2(_11423_),
    .B1(_11306_),
    .B2(_11424_),
    .X(_03506_));
 sky130_fd_sc_hd__a22o_2 _14665_ (.A1(\cpuregs[7][1] ),
    .A2(_11412_),
    .B1(_11307_),
    .B2(_11415_),
    .X(_03505_));
 sky130_fd_sc_hd__a22o_2 _14666_ (.A1(\cpuregs[7][0] ),
    .A2(_11412_),
    .B1(_11308_),
    .B2(_11415_),
    .X(_03504_));
 sky130_vsdinv _14667_ (.A(instr_setq),
    .Y(_11425_));
 sky130_fd_sc_hd__and3_2 _14668_ (.A(_10603_),
    .B(_10606_),
    .C(_00302_),
    .X(_11426_));
 sky130_fd_sc_hd__a2111o_2 _14669_ (.A1(_11425_),
    .A2(_10614_),
    .B1(_10481_),
    .C1(_00331_),
    .D1(_11426_),
    .X(_11427_));
 sky130_fd_sc_hd__mux2_2 _14670_ (.A0(_12943_),
    .A1(\latched_rd[4] ),
    .S(_11427_),
    .X(_03503_));
 sky130_fd_sc_hd__or3_2 _14671_ (.A(\latched_rd[4] ),
    .B(_11309_),
    .C(_11253_),
    .X(_11428_));
 sky130_fd_sc_hd__or2_2 _14672_ (.A(_11381_),
    .B(_11428_),
    .X(_11429_));
 sky130_fd_sc_hd__buf_1 _14673_ (.A(_11429_),
    .X(_11430_));
 sky130_fd_sc_hd__buf_1 _14674_ (.A(_11430_),
    .X(_11431_));
 sky130_vsdinv _14675_ (.A(_11429_),
    .Y(_11432_));
 sky130_fd_sc_hd__buf_1 _14676_ (.A(_11432_),
    .X(_11433_));
 sky130_fd_sc_hd__buf_1 _14677_ (.A(_11433_),
    .X(_11434_));
 sky130_fd_sc_hd__a22o_2 _14678_ (.A1(\cpuregs[15][31] ),
    .A2(_11431_),
    .B1(_11266_),
    .B2(_11434_),
    .X(_03502_));
 sky130_fd_sc_hd__a22o_2 _14679_ (.A1(\cpuregs[15][30] ),
    .A2(_11431_),
    .B1(_11270_),
    .B2(_11434_),
    .X(_03501_));
 sky130_fd_sc_hd__a22o_2 _14680_ (.A1(\cpuregs[15][29] ),
    .A2(_11431_),
    .B1(_11271_),
    .B2(_11434_),
    .X(_03500_));
 sky130_fd_sc_hd__a22o_2 _14681_ (.A1(\cpuregs[15][28] ),
    .A2(_11431_),
    .B1(_11272_),
    .B2(_11434_),
    .X(_03499_));
 sky130_fd_sc_hd__a22o_2 _14682_ (.A1(\cpuregs[15][27] ),
    .A2(_11431_),
    .B1(_11273_),
    .B2(_11434_),
    .X(_03498_));
 sky130_fd_sc_hd__a22o_2 _14683_ (.A1(\cpuregs[15][26] ),
    .A2(_11431_),
    .B1(_11274_),
    .B2(_11434_),
    .X(_03497_));
 sky130_fd_sc_hd__buf_1 _14684_ (.A(_11430_),
    .X(_11435_));
 sky130_fd_sc_hd__buf_1 _14685_ (.A(_11433_),
    .X(_11436_));
 sky130_fd_sc_hd__a22o_2 _14686_ (.A1(\cpuregs[15][25] ),
    .A2(_11435_),
    .B1(_11276_),
    .B2(_11436_),
    .X(_03496_));
 sky130_fd_sc_hd__a22o_2 _14687_ (.A1(\cpuregs[15][24] ),
    .A2(_11435_),
    .B1(_11278_),
    .B2(_11436_),
    .X(_03495_));
 sky130_fd_sc_hd__a22o_2 _14688_ (.A1(\cpuregs[15][23] ),
    .A2(_11435_),
    .B1(_11279_),
    .B2(_11436_),
    .X(_03494_));
 sky130_fd_sc_hd__a22o_2 _14689_ (.A1(\cpuregs[15][22] ),
    .A2(_11435_),
    .B1(_11280_),
    .B2(_11436_),
    .X(_03493_));
 sky130_fd_sc_hd__a22o_2 _14690_ (.A1(\cpuregs[15][21] ),
    .A2(_11435_),
    .B1(_11281_),
    .B2(_11436_),
    .X(_03492_));
 sky130_fd_sc_hd__a22o_2 _14691_ (.A1(\cpuregs[15][20] ),
    .A2(_11435_),
    .B1(_11282_),
    .B2(_11436_),
    .X(_03491_));
 sky130_fd_sc_hd__buf_1 _14692_ (.A(_11430_),
    .X(_11437_));
 sky130_fd_sc_hd__buf_1 _14693_ (.A(_11433_),
    .X(_11438_));
 sky130_fd_sc_hd__a22o_2 _14694_ (.A1(\cpuregs[15][19] ),
    .A2(_11437_),
    .B1(_11284_),
    .B2(_11438_),
    .X(_03490_));
 sky130_fd_sc_hd__a22o_2 _14695_ (.A1(\cpuregs[15][18] ),
    .A2(_11437_),
    .B1(_11286_),
    .B2(_11438_),
    .X(_03489_));
 sky130_fd_sc_hd__a22o_2 _14696_ (.A1(\cpuregs[15][17] ),
    .A2(_11437_),
    .B1(_11287_),
    .B2(_11438_),
    .X(_03488_));
 sky130_fd_sc_hd__a22o_2 _14697_ (.A1(\cpuregs[15][16] ),
    .A2(_11437_),
    .B1(_11288_),
    .B2(_11438_),
    .X(_03487_));
 sky130_fd_sc_hd__a22o_2 _14698_ (.A1(\cpuregs[15][15] ),
    .A2(_11437_),
    .B1(_11289_),
    .B2(_11438_),
    .X(_03486_));
 sky130_fd_sc_hd__a22o_2 _14699_ (.A1(\cpuregs[15][14] ),
    .A2(_11437_),
    .B1(_11290_),
    .B2(_11438_),
    .X(_03485_));
 sky130_fd_sc_hd__buf_1 _14700_ (.A(_11430_),
    .X(_11439_));
 sky130_fd_sc_hd__buf_1 _14701_ (.A(_11433_),
    .X(_11440_));
 sky130_fd_sc_hd__a22o_2 _14702_ (.A1(\cpuregs[15][13] ),
    .A2(_11439_),
    .B1(_11292_),
    .B2(_11440_),
    .X(_03484_));
 sky130_fd_sc_hd__a22o_2 _14703_ (.A1(\cpuregs[15][12] ),
    .A2(_11439_),
    .B1(_11294_),
    .B2(_11440_),
    .X(_03483_));
 sky130_fd_sc_hd__a22o_2 _14704_ (.A1(\cpuregs[15][11] ),
    .A2(_11439_),
    .B1(_11295_),
    .B2(_11440_),
    .X(_03482_));
 sky130_fd_sc_hd__a22o_2 _14705_ (.A1(\cpuregs[15][10] ),
    .A2(_11439_),
    .B1(_11296_),
    .B2(_11440_),
    .X(_03481_));
 sky130_fd_sc_hd__a22o_2 _14706_ (.A1(\cpuregs[15][9] ),
    .A2(_11439_),
    .B1(_11297_),
    .B2(_11440_),
    .X(_03480_));
 sky130_fd_sc_hd__a22o_2 _14707_ (.A1(\cpuregs[15][8] ),
    .A2(_11439_),
    .B1(_11298_),
    .B2(_11440_),
    .X(_03479_));
 sky130_fd_sc_hd__buf_1 _14708_ (.A(_11429_),
    .X(_11441_));
 sky130_fd_sc_hd__buf_1 _14709_ (.A(_11432_),
    .X(_11442_));
 sky130_fd_sc_hd__a22o_2 _14710_ (.A1(\cpuregs[15][7] ),
    .A2(_11441_),
    .B1(_11300_),
    .B2(_11442_),
    .X(_03478_));
 sky130_fd_sc_hd__a22o_2 _14711_ (.A1(\cpuregs[15][6] ),
    .A2(_11441_),
    .B1(_11302_),
    .B2(_11442_),
    .X(_03477_));
 sky130_fd_sc_hd__a22o_2 _14712_ (.A1(\cpuregs[15][5] ),
    .A2(_11441_),
    .B1(_11303_),
    .B2(_11442_),
    .X(_03476_));
 sky130_fd_sc_hd__a22o_2 _14713_ (.A1(\cpuregs[15][4] ),
    .A2(_11441_),
    .B1(_11304_),
    .B2(_11442_),
    .X(_03475_));
 sky130_fd_sc_hd__a22o_2 _14714_ (.A1(\cpuregs[15][3] ),
    .A2(_11441_),
    .B1(_11305_),
    .B2(_11442_),
    .X(_03474_));
 sky130_fd_sc_hd__a22o_2 _14715_ (.A1(\cpuregs[15][2] ),
    .A2(_11441_),
    .B1(_11306_),
    .B2(_11442_),
    .X(_03473_));
 sky130_fd_sc_hd__a22o_2 _14716_ (.A1(\cpuregs[15][1] ),
    .A2(_11430_),
    .B1(_11307_),
    .B2(_11433_),
    .X(_03472_));
 sky130_fd_sc_hd__a22o_2 _14717_ (.A1(\cpuregs[15][0] ),
    .A2(_11430_),
    .B1(_11308_),
    .B2(_11433_),
    .X(_03471_));
 sky130_fd_sc_hd__or2_2 _14718_ (.A(_11311_),
    .B(_11381_),
    .X(_11443_));
 sky130_fd_sc_hd__buf_1 _14719_ (.A(_11443_),
    .X(_11444_));
 sky130_fd_sc_hd__buf_1 _14720_ (.A(_11444_),
    .X(_11445_));
 sky130_fd_sc_hd__buf_1 _14721_ (.A(\cpuregs_wrdata[31] ),
    .X(_11446_));
 sky130_vsdinv _14722_ (.A(_11443_),
    .Y(_11447_));
 sky130_fd_sc_hd__buf_1 _14723_ (.A(_11447_),
    .X(_11448_));
 sky130_fd_sc_hd__buf_1 _14724_ (.A(_11448_),
    .X(_11449_));
 sky130_fd_sc_hd__a22o_2 _14725_ (.A1(\cpuregs[11][31] ),
    .A2(_11445_),
    .B1(_11446_),
    .B2(_11449_),
    .X(_03470_));
 sky130_fd_sc_hd__buf_1 _14726_ (.A(\cpuregs_wrdata[30] ),
    .X(_11450_));
 sky130_fd_sc_hd__a22o_2 _14727_ (.A1(\cpuregs[11][30] ),
    .A2(_11445_),
    .B1(_11450_),
    .B2(_11449_),
    .X(_03469_));
 sky130_fd_sc_hd__buf_1 _14728_ (.A(\cpuregs_wrdata[29] ),
    .X(_11451_));
 sky130_fd_sc_hd__a22o_2 _14729_ (.A1(\cpuregs[11][29] ),
    .A2(_11445_),
    .B1(_11451_),
    .B2(_11449_),
    .X(_03468_));
 sky130_fd_sc_hd__buf_1 _14730_ (.A(\cpuregs_wrdata[28] ),
    .X(_11452_));
 sky130_fd_sc_hd__a22o_2 _14731_ (.A1(\cpuregs[11][28] ),
    .A2(_11445_),
    .B1(_11452_),
    .B2(_11449_),
    .X(_03467_));
 sky130_fd_sc_hd__buf_1 _14732_ (.A(\cpuregs_wrdata[27] ),
    .X(_11453_));
 sky130_fd_sc_hd__a22o_2 _14733_ (.A1(\cpuregs[11][27] ),
    .A2(_11445_),
    .B1(_11453_),
    .B2(_11449_),
    .X(_03466_));
 sky130_fd_sc_hd__buf_1 _14734_ (.A(\cpuregs_wrdata[26] ),
    .X(_11454_));
 sky130_fd_sc_hd__a22o_2 _14735_ (.A1(\cpuregs[11][26] ),
    .A2(_11445_),
    .B1(_11454_),
    .B2(_11449_),
    .X(_03465_));
 sky130_fd_sc_hd__buf_1 _14736_ (.A(_11444_),
    .X(_11455_));
 sky130_fd_sc_hd__buf_1 _14737_ (.A(\cpuregs_wrdata[25] ),
    .X(_11456_));
 sky130_fd_sc_hd__buf_1 _14738_ (.A(_11448_),
    .X(_11457_));
 sky130_fd_sc_hd__a22o_2 _14739_ (.A1(\cpuregs[11][25] ),
    .A2(_11455_),
    .B1(_11456_),
    .B2(_11457_),
    .X(_03464_));
 sky130_fd_sc_hd__buf_1 _14740_ (.A(\cpuregs_wrdata[24] ),
    .X(_11458_));
 sky130_fd_sc_hd__a22o_2 _14741_ (.A1(\cpuregs[11][24] ),
    .A2(_11455_),
    .B1(_11458_),
    .B2(_11457_),
    .X(_03463_));
 sky130_fd_sc_hd__buf_1 _14742_ (.A(\cpuregs_wrdata[23] ),
    .X(_11459_));
 sky130_fd_sc_hd__a22o_2 _14743_ (.A1(\cpuregs[11][23] ),
    .A2(_11455_),
    .B1(_11459_),
    .B2(_11457_),
    .X(_03462_));
 sky130_fd_sc_hd__buf_1 _14744_ (.A(\cpuregs_wrdata[22] ),
    .X(_11460_));
 sky130_fd_sc_hd__a22o_2 _14745_ (.A1(\cpuregs[11][22] ),
    .A2(_11455_),
    .B1(_11460_),
    .B2(_11457_),
    .X(_03461_));
 sky130_fd_sc_hd__buf_1 _14746_ (.A(\cpuregs_wrdata[21] ),
    .X(_11461_));
 sky130_fd_sc_hd__a22o_2 _14747_ (.A1(\cpuregs[11][21] ),
    .A2(_11455_),
    .B1(_11461_),
    .B2(_11457_),
    .X(_03460_));
 sky130_fd_sc_hd__buf_1 _14748_ (.A(\cpuregs_wrdata[20] ),
    .X(_11462_));
 sky130_fd_sc_hd__a22o_2 _14749_ (.A1(\cpuregs[11][20] ),
    .A2(_11455_),
    .B1(_11462_),
    .B2(_11457_),
    .X(_03459_));
 sky130_fd_sc_hd__buf_1 _14750_ (.A(_11444_),
    .X(_11463_));
 sky130_fd_sc_hd__buf_1 _14751_ (.A(\cpuregs_wrdata[19] ),
    .X(_11464_));
 sky130_fd_sc_hd__buf_1 _14752_ (.A(_11448_),
    .X(_11465_));
 sky130_fd_sc_hd__a22o_2 _14753_ (.A1(\cpuregs[11][19] ),
    .A2(_11463_),
    .B1(_11464_),
    .B2(_11465_),
    .X(_03458_));
 sky130_fd_sc_hd__buf_1 _14754_ (.A(\cpuregs_wrdata[18] ),
    .X(_11466_));
 sky130_fd_sc_hd__a22o_2 _14755_ (.A1(\cpuregs[11][18] ),
    .A2(_11463_),
    .B1(_11466_),
    .B2(_11465_),
    .X(_03457_));
 sky130_fd_sc_hd__buf_1 _14756_ (.A(\cpuregs_wrdata[17] ),
    .X(_11467_));
 sky130_fd_sc_hd__a22o_2 _14757_ (.A1(\cpuregs[11][17] ),
    .A2(_11463_),
    .B1(_11467_),
    .B2(_11465_),
    .X(_03456_));
 sky130_fd_sc_hd__buf_1 _14758_ (.A(\cpuregs_wrdata[16] ),
    .X(_11468_));
 sky130_fd_sc_hd__a22o_2 _14759_ (.A1(\cpuregs[11][16] ),
    .A2(_11463_),
    .B1(_11468_),
    .B2(_11465_),
    .X(_03455_));
 sky130_fd_sc_hd__buf_1 _14760_ (.A(\cpuregs_wrdata[15] ),
    .X(_11469_));
 sky130_fd_sc_hd__a22o_2 _14761_ (.A1(\cpuregs[11][15] ),
    .A2(_11463_),
    .B1(_11469_),
    .B2(_11465_),
    .X(_03454_));
 sky130_fd_sc_hd__buf_1 _14762_ (.A(\cpuregs_wrdata[14] ),
    .X(_11470_));
 sky130_fd_sc_hd__a22o_2 _14763_ (.A1(\cpuregs[11][14] ),
    .A2(_11463_),
    .B1(_11470_),
    .B2(_11465_),
    .X(_03453_));
 sky130_fd_sc_hd__buf_1 _14764_ (.A(_11444_),
    .X(_11471_));
 sky130_fd_sc_hd__buf_1 _14765_ (.A(\cpuregs_wrdata[13] ),
    .X(_11472_));
 sky130_fd_sc_hd__buf_1 _14766_ (.A(_11448_),
    .X(_11473_));
 sky130_fd_sc_hd__a22o_2 _14767_ (.A1(\cpuregs[11][13] ),
    .A2(_11471_),
    .B1(_11472_),
    .B2(_11473_),
    .X(_03452_));
 sky130_fd_sc_hd__buf_1 _14768_ (.A(\cpuregs_wrdata[12] ),
    .X(_11474_));
 sky130_fd_sc_hd__a22o_2 _14769_ (.A1(\cpuregs[11][12] ),
    .A2(_11471_),
    .B1(_11474_),
    .B2(_11473_),
    .X(_03451_));
 sky130_fd_sc_hd__buf_1 _14770_ (.A(\cpuregs_wrdata[11] ),
    .X(_11475_));
 sky130_fd_sc_hd__a22o_2 _14771_ (.A1(\cpuregs[11][11] ),
    .A2(_11471_),
    .B1(_11475_),
    .B2(_11473_),
    .X(_03450_));
 sky130_fd_sc_hd__buf_1 _14772_ (.A(\cpuregs_wrdata[10] ),
    .X(_11476_));
 sky130_fd_sc_hd__a22o_2 _14773_ (.A1(\cpuregs[11][10] ),
    .A2(_11471_),
    .B1(_11476_),
    .B2(_11473_),
    .X(_03449_));
 sky130_fd_sc_hd__buf_1 _14774_ (.A(\cpuregs_wrdata[9] ),
    .X(_11477_));
 sky130_fd_sc_hd__a22o_2 _14775_ (.A1(\cpuregs[11][9] ),
    .A2(_11471_),
    .B1(_11477_),
    .B2(_11473_),
    .X(_03448_));
 sky130_fd_sc_hd__buf_1 _14776_ (.A(\cpuregs_wrdata[8] ),
    .X(_11478_));
 sky130_fd_sc_hd__a22o_2 _14777_ (.A1(\cpuregs[11][8] ),
    .A2(_11471_),
    .B1(_11478_),
    .B2(_11473_),
    .X(_03447_));
 sky130_fd_sc_hd__buf_1 _14778_ (.A(_11443_),
    .X(_11479_));
 sky130_fd_sc_hd__buf_1 _14779_ (.A(\cpuregs_wrdata[7] ),
    .X(_11480_));
 sky130_fd_sc_hd__buf_1 _14780_ (.A(_11447_),
    .X(_11481_));
 sky130_fd_sc_hd__a22o_2 _14781_ (.A1(\cpuregs[11][7] ),
    .A2(_11479_),
    .B1(_11480_),
    .B2(_11481_),
    .X(_03446_));
 sky130_fd_sc_hd__buf_1 _14782_ (.A(\cpuregs_wrdata[6] ),
    .X(_11482_));
 sky130_fd_sc_hd__a22o_2 _14783_ (.A1(\cpuregs[11][6] ),
    .A2(_11479_),
    .B1(_11482_),
    .B2(_11481_),
    .X(_03445_));
 sky130_fd_sc_hd__buf_1 _14784_ (.A(\cpuregs_wrdata[5] ),
    .X(_11483_));
 sky130_fd_sc_hd__a22o_2 _14785_ (.A1(\cpuregs[11][5] ),
    .A2(_11479_),
    .B1(_11483_),
    .B2(_11481_),
    .X(_03444_));
 sky130_fd_sc_hd__buf_1 _14786_ (.A(\cpuregs_wrdata[4] ),
    .X(_11484_));
 sky130_fd_sc_hd__a22o_2 _14787_ (.A1(\cpuregs[11][4] ),
    .A2(_11479_),
    .B1(_11484_),
    .B2(_11481_),
    .X(_03443_));
 sky130_fd_sc_hd__buf_1 _14788_ (.A(\cpuregs_wrdata[3] ),
    .X(_11485_));
 sky130_fd_sc_hd__a22o_2 _14789_ (.A1(\cpuregs[11][3] ),
    .A2(_11479_),
    .B1(_11485_),
    .B2(_11481_),
    .X(_03442_));
 sky130_fd_sc_hd__buf_1 _14790_ (.A(\cpuregs_wrdata[2] ),
    .X(_11486_));
 sky130_fd_sc_hd__a22o_2 _14791_ (.A1(\cpuregs[11][2] ),
    .A2(_11479_),
    .B1(_11486_),
    .B2(_11481_),
    .X(_03441_));
 sky130_fd_sc_hd__buf_1 _14792_ (.A(\cpuregs_wrdata[1] ),
    .X(_11487_));
 sky130_fd_sc_hd__a22o_2 _14793_ (.A1(\cpuregs[11][1] ),
    .A2(_11444_),
    .B1(_11487_),
    .B2(_11448_),
    .X(_03440_));
 sky130_fd_sc_hd__buf_1 _14794_ (.A(\cpuregs_wrdata[0] ),
    .X(_11488_));
 sky130_fd_sc_hd__a22o_2 _14795_ (.A1(\cpuregs[11][0] ),
    .A2(_11444_),
    .B1(_11488_),
    .B2(_11448_),
    .X(_03439_));
 sky130_fd_sc_hd__or2_2 _14796_ (.A(_11258_),
    .B(_11381_),
    .X(_11489_));
 sky130_fd_sc_hd__buf_1 _14797_ (.A(_11489_),
    .X(_11490_));
 sky130_fd_sc_hd__buf_1 _14798_ (.A(_11490_),
    .X(_11491_));
 sky130_vsdinv _14799_ (.A(_11489_),
    .Y(_11492_));
 sky130_fd_sc_hd__buf_1 _14800_ (.A(_11492_),
    .X(_11493_));
 sky130_fd_sc_hd__buf_1 _14801_ (.A(_11493_),
    .X(_11494_));
 sky130_fd_sc_hd__a22o_2 _14802_ (.A1(\cpuregs[3][31] ),
    .A2(_11491_),
    .B1(_11446_),
    .B2(_11494_),
    .X(_03438_));
 sky130_fd_sc_hd__a22o_2 _14803_ (.A1(\cpuregs[3][30] ),
    .A2(_11491_),
    .B1(_11450_),
    .B2(_11494_),
    .X(_03437_));
 sky130_fd_sc_hd__a22o_2 _14804_ (.A1(\cpuregs[3][29] ),
    .A2(_11491_),
    .B1(_11451_),
    .B2(_11494_),
    .X(_03436_));
 sky130_fd_sc_hd__a22o_2 _14805_ (.A1(\cpuregs[3][28] ),
    .A2(_11491_),
    .B1(_11452_),
    .B2(_11494_),
    .X(_03435_));
 sky130_fd_sc_hd__a22o_2 _14806_ (.A1(\cpuregs[3][27] ),
    .A2(_11491_),
    .B1(_11453_),
    .B2(_11494_),
    .X(_03434_));
 sky130_fd_sc_hd__a22o_2 _14807_ (.A1(\cpuregs[3][26] ),
    .A2(_11491_),
    .B1(_11454_),
    .B2(_11494_),
    .X(_03433_));
 sky130_fd_sc_hd__buf_1 _14808_ (.A(_11490_),
    .X(_11495_));
 sky130_fd_sc_hd__buf_1 _14809_ (.A(_11493_),
    .X(_11496_));
 sky130_fd_sc_hd__a22o_2 _14810_ (.A1(\cpuregs[3][25] ),
    .A2(_11495_),
    .B1(_11456_),
    .B2(_11496_),
    .X(_03432_));
 sky130_fd_sc_hd__a22o_2 _14811_ (.A1(\cpuregs[3][24] ),
    .A2(_11495_),
    .B1(_11458_),
    .B2(_11496_),
    .X(_03431_));
 sky130_fd_sc_hd__a22o_2 _14812_ (.A1(\cpuregs[3][23] ),
    .A2(_11495_),
    .B1(_11459_),
    .B2(_11496_),
    .X(_03430_));
 sky130_fd_sc_hd__a22o_2 _14813_ (.A1(\cpuregs[3][22] ),
    .A2(_11495_),
    .B1(_11460_),
    .B2(_11496_),
    .X(_03429_));
 sky130_fd_sc_hd__a22o_2 _14814_ (.A1(\cpuregs[3][21] ),
    .A2(_11495_),
    .B1(_11461_),
    .B2(_11496_),
    .X(_03428_));
 sky130_fd_sc_hd__a22o_2 _14815_ (.A1(\cpuregs[3][20] ),
    .A2(_11495_),
    .B1(_11462_),
    .B2(_11496_),
    .X(_03427_));
 sky130_fd_sc_hd__buf_1 _14816_ (.A(_11490_),
    .X(_11497_));
 sky130_fd_sc_hd__buf_1 _14817_ (.A(_11493_),
    .X(_11498_));
 sky130_fd_sc_hd__a22o_2 _14818_ (.A1(\cpuregs[3][19] ),
    .A2(_11497_),
    .B1(_11464_),
    .B2(_11498_),
    .X(_03426_));
 sky130_fd_sc_hd__a22o_2 _14819_ (.A1(\cpuregs[3][18] ),
    .A2(_11497_),
    .B1(_11466_),
    .B2(_11498_),
    .X(_03425_));
 sky130_fd_sc_hd__a22o_2 _14820_ (.A1(\cpuregs[3][17] ),
    .A2(_11497_),
    .B1(_11467_),
    .B2(_11498_),
    .X(_03424_));
 sky130_fd_sc_hd__a22o_2 _14821_ (.A1(\cpuregs[3][16] ),
    .A2(_11497_),
    .B1(_11468_),
    .B2(_11498_),
    .X(_03423_));
 sky130_fd_sc_hd__a22o_2 _14822_ (.A1(\cpuregs[3][15] ),
    .A2(_11497_),
    .B1(_11469_),
    .B2(_11498_),
    .X(_03422_));
 sky130_fd_sc_hd__a22o_2 _14823_ (.A1(\cpuregs[3][14] ),
    .A2(_11497_),
    .B1(_11470_),
    .B2(_11498_),
    .X(_03421_));
 sky130_fd_sc_hd__buf_1 _14824_ (.A(_11490_),
    .X(_11499_));
 sky130_fd_sc_hd__buf_1 _14825_ (.A(_11493_),
    .X(_11500_));
 sky130_fd_sc_hd__a22o_2 _14826_ (.A1(\cpuregs[3][13] ),
    .A2(_11499_),
    .B1(_11472_),
    .B2(_11500_),
    .X(_03420_));
 sky130_fd_sc_hd__a22o_2 _14827_ (.A1(\cpuregs[3][12] ),
    .A2(_11499_),
    .B1(_11474_),
    .B2(_11500_),
    .X(_03419_));
 sky130_fd_sc_hd__a22o_2 _14828_ (.A1(\cpuregs[3][11] ),
    .A2(_11499_),
    .B1(_11475_),
    .B2(_11500_),
    .X(_03418_));
 sky130_fd_sc_hd__a22o_2 _14829_ (.A1(\cpuregs[3][10] ),
    .A2(_11499_),
    .B1(_11476_),
    .B2(_11500_),
    .X(_03417_));
 sky130_fd_sc_hd__a22o_2 _14830_ (.A1(\cpuregs[3][9] ),
    .A2(_11499_),
    .B1(_11477_),
    .B2(_11500_),
    .X(_03416_));
 sky130_fd_sc_hd__a22o_2 _14831_ (.A1(\cpuregs[3][8] ),
    .A2(_11499_),
    .B1(_11478_),
    .B2(_11500_),
    .X(_03415_));
 sky130_fd_sc_hd__buf_1 _14832_ (.A(_11489_),
    .X(_11501_));
 sky130_fd_sc_hd__buf_1 _14833_ (.A(_11492_),
    .X(_11502_));
 sky130_fd_sc_hd__a22o_2 _14834_ (.A1(\cpuregs[3][7] ),
    .A2(_11501_),
    .B1(_11480_),
    .B2(_11502_),
    .X(_03414_));
 sky130_fd_sc_hd__a22o_2 _14835_ (.A1(\cpuregs[3][6] ),
    .A2(_11501_),
    .B1(_11482_),
    .B2(_11502_),
    .X(_03413_));
 sky130_fd_sc_hd__a22o_2 _14836_ (.A1(\cpuregs[3][5] ),
    .A2(_11501_),
    .B1(_11483_),
    .B2(_11502_),
    .X(_03412_));
 sky130_fd_sc_hd__a22o_2 _14837_ (.A1(\cpuregs[3][4] ),
    .A2(_11501_),
    .B1(_11484_),
    .B2(_11502_),
    .X(_03411_));
 sky130_fd_sc_hd__a22o_2 _14838_ (.A1(\cpuregs[3][3] ),
    .A2(_11501_),
    .B1(_11485_),
    .B2(_11502_),
    .X(_03410_));
 sky130_fd_sc_hd__a22o_2 _14839_ (.A1(\cpuregs[3][2] ),
    .A2(_11501_),
    .B1(_11486_),
    .B2(_11502_),
    .X(_03409_));
 sky130_fd_sc_hd__a22o_2 _14840_ (.A1(\cpuregs[3][1] ),
    .A2(_11490_),
    .B1(_11487_),
    .B2(_11493_),
    .X(_03408_));
 sky130_fd_sc_hd__a22o_2 _14841_ (.A1(\cpuregs[3][0] ),
    .A2(_11490_),
    .B1(_11488_),
    .B2(_11493_),
    .X(_03407_));
 sky130_fd_sc_hd__or2_2 _14842_ (.A(_11258_),
    .B(_11313_),
    .X(_11503_));
 sky130_fd_sc_hd__buf_1 _14843_ (.A(_11503_),
    .X(_11504_));
 sky130_fd_sc_hd__buf_1 _14844_ (.A(_11504_),
    .X(_11505_));
 sky130_vsdinv _14845_ (.A(_11503_),
    .Y(_11506_));
 sky130_fd_sc_hd__buf_1 _14846_ (.A(_11506_),
    .X(_11507_));
 sky130_fd_sc_hd__buf_1 _14847_ (.A(_11507_),
    .X(_11508_));
 sky130_fd_sc_hd__a22o_2 _14848_ (.A1(\cpuregs[1][31] ),
    .A2(_11505_),
    .B1(_11446_),
    .B2(_11508_),
    .X(_03406_));
 sky130_fd_sc_hd__a22o_2 _14849_ (.A1(\cpuregs[1][30] ),
    .A2(_11505_),
    .B1(_11450_),
    .B2(_11508_),
    .X(_03405_));
 sky130_fd_sc_hd__a22o_2 _14850_ (.A1(\cpuregs[1][29] ),
    .A2(_11505_),
    .B1(_11451_),
    .B2(_11508_),
    .X(_03404_));
 sky130_fd_sc_hd__a22o_2 _14851_ (.A1(\cpuregs[1][28] ),
    .A2(_11505_),
    .B1(_11452_),
    .B2(_11508_),
    .X(_03403_));
 sky130_fd_sc_hd__a22o_2 _14852_ (.A1(\cpuregs[1][27] ),
    .A2(_11505_),
    .B1(_11453_),
    .B2(_11508_),
    .X(_03402_));
 sky130_fd_sc_hd__a22o_2 _14853_ (.A1(\cpuregs[1][26] ),
    .A2(_11505_),
    .B1(_11454_),
    .B2(_11508_),
    .X(_03401_));
 sky130_fd_sc_hd__buf_1 _14854_ (.A(_11504_),
    .X(_11509_));
 sky130_fd_sc_hd__buf_1 _14855_ (.A(_11507_),
    .X(_11510_));
 sky130_fd_sc_hd__a22o_2 _14856_ (.A1(\cpuregs[1][25] ),
    .A2(_11509_),
    .B1(_11456_),
    .B2(_11510_),
    .X(_03400_));
 sky130_fd_sc_hd__a22o_2 _14857_ (.A1(\cpuregs[1][24] ),
    .A2(_11509_),
    .B1(_11458_),
    .B2(_11510_),
    .X(_03399_));
 sky130_fd_sc_hd__a22o_2 _14858_ (.A1(\cpuregs[1][23] ),
    .A2(_11509_),
    .B1(_11459_),
    .B2(_11510_),
    .X(_03398_));
 sky130_fd_sc_hd__a22o_2 _14859_ (.A1(\cpuregs[1][22] ),
    .A2(_11509_),
    .B1(_11460_),
    .B2(_11510_),
    .X(_03397_));
 sky130_fd_sc_hd__a22o_2 _14860_ (.A1(\cpuregs[1][21] ),
    .A2(_11509_),
    .B1(_11461_),
    .B2(_11510_),
    .X(_03396_));
 sky130_fd_sc_hd__a22o_2 _14861_ (.A1(\cpuregs[1][20] ),
    .A2(_11509_),
    .B1(_11462_),
    .B2(_11510_),
    .X(_03395_));
 sky130_fd_sc_hd__buf_1 _14862_ (.A(_11504_),
    .X(_11511_));
 sky130_fd_sc_hd__buf_1 _14863_ (.A(_11507_),
    .X(_11512_));
 sky130_fd_sc_hd__a22o_2 _14864_ (.A1(\cpuregs[1][19] ),
    .A2(_11511_),
    .B1(_11464_),
    .B2(_11512_),
    .X(_03394_));
 sky130_fd_sc_hd__a22o_2 _14865_ (.A1(\cpuregs[1][18] ),
    .A2(_11511_),
    .B1(_11466_),
    .B2(_11512_),
    .X(_03393_));
 sky130_fd_sc_hd__a22o_2 _14866_ (.A1(\cpuregs[1][17] ),
    .A2(_11511_),
    .B1(_11467_),
    .B2(_11512_),
    .X(_03392_));
 sky130_fd_sc_hd__a22o_2 _14867_ (.A1(\cpuregs[1][16] ),
    .A2(_11511_),
    .B1(_11468_),
    .B2(_11512_),
    .X(_03391_));
 sky130_fd_sc_hd__a22o_2 _14868_ (.A1(\cpuregs[1][15] ),
    .A2(_11511_),
    .B1(_11469_),
    .B2(_11512_),
    .X(_03390_));
 sky130_fd_sc_hd__a22o_2 _14869_ (.A1(\cpuregs[1][14] ),
    .A2(_11511_),
    .B1(_11470_),
    .B2(_11512_),
    .X(_03389_));
 sky130_fd_sc_hd__buf_1 _14870_ (.A(_11504_),
    .X(_11513_));
 sky130_fd_sc_hd__buf_1 _14871_ (.A(_11507_),
    .X(_11514_));
 sky130_fd_sc_hd__a22o_2 _14872_ (.A1(\cpuregs[1][13] ),
    .A2(_11513_),
    .B1(_11472_),
    .B2(_11514_),
    .X(_03388_));
 sky130_fd_sc_hd__a22o_2 _14873_ (.A1(\cpuregs[1][12] ),
    .A2(_11513_),
    .B1(_11474_),
    .B2(_11514_),
    .X(_03387_));
 sky130_fd_sc_hd__a22o_2 _14874_ (.A1(\cpuregs[1][11] ),
    .A2(_11513_),
    .B1(_11475_),
    .B2(_11514_),
    .X(_03386_));
 sky130_fd_sc_hd__a22o_2 _14875_ (.A1(\cpuregs[1][10] ),
    .A2(_11513_),
    .B1(_11476_),
    .B2(_11514_),
    .X(_03385_));
 sky130_fd_sc_hd__a22o_2 _14876_ (.A1(\cpuregs[1][9] ),
    .A2(_11513_),
    .B1(_11477_),
    .B2(_11514_),
    .X(_03384_));
 sky130_fd_sc_hd__a22o_2 _14877_ (.A1(\cpuregs[1][8] ),
    .A2(_11513_),
    .B1(_11478_),
    .B2(_11514_),
    .X(_03383_));
 sky130_fd_sc_hd__buf_1 _14878_ (.A(_11503_),
    .X(_11515_));
 sky130_fd_sc_hd__buf_1 _14879_ (.A(_11506_),
    .X(_11516_));
 sky130_fd_sc_hd__a22o_2 _14880_ (.A1(\cpuregs[1][7] ),
    .A2(_11515_),
    .B1(_11480_),
    .B2(_11516_),
    .X(_03382_));
 sky130_fd_sc_hd__a22o_2 _14881_ (.A1(\cpuregs[1][6] ),
    .A2(_11515_),
    .B1(_11482_),
    .B2(_11516_),
    .X(_03381_));
 sky130_fd_sc_hd__a22o_2 _14882_ (.A1(\cpuregs[1][5] ),
    .A2(_11515_),
    .B1(_11483_),
    .B2(_11516_),
    .X(_03380_));
 sky130_fd_sc_hd__a22o_2 _14883_ (.A1(\cpuregs[1][4] ),
    .A2(_11515_),
    .B1(_11484_),
    .B2(_11516_),
    .X(_03379_));
 sky130_fd_sc_hd__a22o_2 _14884_ (.A1(\cpuregs[1][3] ),
    .A2(_11515_),
    .B1(_11485_),
    .B2(_11516_),
    .X(_03378_));
 sky130_fd_sc_hd__a22o_2 _14885_ (.A1(\cpuregs[1][2] ),
    .A2(_11515_),
    .B1(_11486_),
    .B2(_11516_),
    .X(_03377_));
 sky130_fd_sc_hd__a22o_2 _14886_ (.A1(\cpuregs[1][1] ),
    .A2(_11504_),
    .B1(_11487_),
    .B2(_11507_),
    .X(_03376_));
 sky130_fd_sc_hd__a22o_2 _14887_ (.A1(\cpuregs[1][0] ),
    .A2(_11504_),
    .B1(_11488_),
    .B2(_11507_),
    .X(_03375_));
 sky130_fd_sc_hd__or2_2 _14888_ (.A(_11365_),
    .B(_11428_),
    .X(_11517_));
 sky130_fd_sc_hd__buf_1 _14889_ (.A(_11517_),
    .X(_11518_));
 sky130_fd_sc_hd__buf_1 _14890_ (.A(_11518_),
    .X(_11519_));
 sky130_vsdinv _14891_ (.A(_11517_),
    .Y(_11520_));
 sky130_fd_sc_hd__buf_1 _14892_ (.A(_11520_),
    .X(_11521_));
 sky130_fd_sc_hd__buf_1 _14893_ (.A(_11521_),
    .X(_11522_));
 sky130_fd_sc_hd__a22o_2 _14894_ (.A1(\cpuregs[12][31] ),
    .A2(_11519_),
    .B1(_11446_),
    .B2(_11522_),
    .X(_03374_));
 sky130_fd_sc_hd__a22o_2 _14895_ (.A1(\cpuregs[12][30] ),
    .A2(_11519_),
    .B1(_11450_),
    .B2(_11522_),
    .X(_03373_));
 sky130_fd_sc_hd__a22o_2 _14896_ (.A1(\cpuregs[12][29] ),
    .A2(_11519_),
    .B1(_11451_),
    .B2(_11522_),
    .X(_03372_));
 sky130_fd_sc_hd__a22o_2 _14897_ (.A1(\cpuregs[12][28] ),
    .A2(_11519_),
    .B1(_11452_),
    .B2(_11522_),
    .X(_03371_));
 sky130_fd_sc_hd__a22o_2 _14898_ (.A1(\cpuregs[12][27] ),
    .A2(_11519_),
    .B1(_11453_),
    .B2(_11522_),
    .X(_03370_));
 sky130_fd_sc_hd__a22o_2 _14899_ (.A1(\cpuregs[12][26] ),
    .A2(_11519_),
    .B1(_11454_),
    .B2(_11522_),
    .X(_03369_));
 sky130_fd_sc_hd__buf_1 _14900_ (.A(_11518_),
    .X(_11523_));
 sky130_fd_sc_hd__buf_1 _14901_ (.A(_11521_),
    .X(_11524_));
 sky130_fd_sc_hd__a22o_2 _14902_ (.A1(\cpuregs[12][25] ),
    .A2(_11523_),
    .B1(_11456_),
    .B2(_11524_),
    .X(_03368_));
 sky130_fd_sc_hd__a22o_2 _14903_ (.A1(\cpuregs[12][24] ),
    .A2(_11523_),
    .B1(_11458_),
    .B2(_11524_),
    .X(_03367_));
 sky130_fd_sc_hd__a22o_2 _14904_ (.A1(\cpuregs[12][23] ),
    .A2(_11523_),
    .B1(_11459_),
    .B2(_11524_),
    .X(_03366_));
 sky130_fd_sc_hd__a22o_2 _14905_ (.A1(\cpuregs[12][22] ),
    .A2(_11523_),
    .B1(_11460_),
    .B2(_11524_),
    .X(_03365_));
 sky130_fd_sc_hd__a22o_2 _14906_ (.A1(\cpuregs[12][21] ),
    .A2(_11523_),
    .B1(_11461_),
    .B2(_11524_),
    .X(_03364_));
 sky130_fd_sc_hd__a22o_2 _14907_ (.A1(\cpuregs[12][20] ),
    .A2(_11523_),
    .B1(_11462_),
    .B2(_11524_),
    .X(_03363_));
 sky130_fd_sc_hd__buf_1 _14908_ (.A(_11518_),
    .X(_11525_));
 sky130_fd_sc_hd__buf_1 _14909_ (.A(_11521_),
    .X(_11526_));
 sky130_fd_sc_hd__a22o_2 _14910_ (.A1(\cpuregs[12][19] ),
    .A2(_11525_),
    .B1(_11464_),
    .B2(_11526_),
    .X(_03362_));
 sky130_fd_sc_hd__a22o_2 _14911_ (.A1(\cpuregs[12][18] ),
    .A2(_11525_),
    .B1(_11466_),
    .B2(_11526_),
    .X(_03361_));
 sky130_fd_sc_hd__a22o_2 _14912_ (.A1(\cpuregs[12][17] ),
    .A2(_11525_),
    .B1(_11467_),
    .B2(_11526_),
    .X(_03360_));
 sky130_fd_sc_hd__a22o_2 _14913_ (.A1(\cpuregs[12][16] ),
    .A2(_11525_),
    .B1(_11468_),
    .B2(_11526_),
    .X(_03359_));
 sky130_fd_sc_hd__a22o_2 _14914_ (.A1(\cpuregs[12][15] ),
    .A2(_11525_),
    .B1(_11469_),
    .B2(_11526_),
    .X(_03358_));
 sky130_fd_sc_hd__a22o_2 _14915_ (.A1(\cpuregs[12][14] ),
    .A2(_11525_),
    .B1(_11470_),
    .B2(_11526_),
    .X(_03357_));
 sky130_fd_sc_hd__buf_1 _14916_ (.A(_11518_),
    .X(_11527_));
 sky130_fd_sc_hd__buf_1 _14917_ (.A(_11521_),
    .X(_11528_));
 sky130_fd_sc_hd__a22o_2 _14918_ (.A1(\cpuregs[12][13] ),
    .A2(_11527_),
    .B1(_11472_),
    .B2(_11528_),
    .X(_03356_));
 sky130_fd_sc_hd__a22o_2 _14919_ (.A1(\cpuregs[12][12] ),
    .A2(_11527_),
    .B1(_11474_),
    .B2(_11528_),
    .X(_03355_));
 sky130_fd_sc_hd__a22o_2 _14920_ (.A1(\cpuregs[12][11] ),
    .A2(_11527_),
    .B1(_11475_),
    .B2(_11528_),
    .X(_03354_));
 sky130_fd_sc_hd__a22o_2 _14921_ (.A1(\cpuregs[12][10] ),
    .A2(_11527_),
    .B1(_11476_),
    .B2(_11528_),
    .X(_03353_));
 sky130_fd_sc_hd__a22o_2 _14922_ (.A1(\cpuregs[12][9] ),
    .A2(_11527_),
    .B1(_11477_),
    .B2(_11528_),
    .X(_03352_));
 sky130_fd_sc_hd__a22o_2 _14923_ (.A1(\cpuregs[12][8] ),
    .A2(_11527_),
    .B1(_11478_),
    .B2(_11528_),
    .X(_03351_));
 sky130_fd_sc_hd__buf_1 _14924_ (.A(_11517_),
    .X(_11529_));
 sky130_fd_sc_hd__buf_1 _14925_ (.A(_11520_),
    .X(_11530_));
 sky130_fd_sc_hd__a22o_2 _14926_ (.A1(\cpuregs[12][7] ),
    .A2(_11529_),
    .B1(_11480_),
    .B2(_11530_),
    .X(_03350_));
 sky130_fd_sc_hd__a22o_2 _14927_ (.A1(\cpuregs[12][6] ),
    .A2(_11529_),
    .B1(_11482_),
    .B2(_11530_),
    .X(_03349_));
 sky130_fd_sc_hd__a22o_2 _14928_ (.A1(\cpuregs[12][5] ),
    .A2(_11529_),
    .B1(_11483_),
    .B2(_11530_),
    .X(_03348_));
 sky130_fd_sc_hd__a22o_2 _14929_ (.A1(\cpuregs[12][4] ),
    .A2(_11529_),
    .B1(_11484_),
    .B2(_11530_),
    .X(_03347_));
 sky130_fd_sc_hd__a22o_2 _14930_ (.A1(\cpuregs[12][3] ),
    .A2(_11529_),
    .B1(_11485_),
    .B2(_11530_),
    .X(_03346_));
 sky130_fd_sc_hd__a22o_2 _14931_ (.A1(\cpuregs[12][2] ),
    .A2(_11529_),
    .B1(_11486_),
    .B2(_11530_),
    .X(_03345_));
 sky130_fd_sc_hd__a22o_2 _14932_ (.A1(\cpuregs[12][1] ),
    .A2(_11518_),
    .B1(_11487_),
    .B2(_11521_),
    .X(_03344_));
 sky130_fd_sc_hd__a22o_2 _14933_ (.A1(\cpuregs[12][0] ),
    .A2(_11518_),
    .B1(_11488_),
    .B2(_11521_),
    .X(_03343_));
 sky130_fd_sc_hd__or3_2 _14934_ (.A(_11310_),
    .B(_11252_),
    .C(_11365_),
    .X(_11531_));
 sky130_fd_sc_hd__buf_1 _14935_ (.A(_11531_),
    .X(_11532_));
 sky130_fd_sc_hd__buf_1 _14936_ (.A(_11532_),
    .X(_11533_));
 sky130_vsdinv _14937_ (.A(_11531_),
    .Y(_11534_));
 sky130_fd_sc_hd__buf_1 _14938_ (.A(_11534_),
    .X(_11535_));
 sky130_fd_sc_hd__buf_1 _14939_ (.A(_11535_),
    .X(_11536_));
 sky130_fd_sc_hd__a22o_2 _14940_ (.A1(\cpuregs[16][31] ),
    .A2(_11533_),
    .B1(_11446_),
    .B2(_11536_),
    .X(_03342_));
 sky130_fd_sc_hd__a22o_2 _14941_ (.A1(\cpuregs[16][30] ),
    .A2(_11533_),
    .B1(_11450_),
    .B2(_11536_),
    .X(_03341_));
 sky130_fd_sc_hd__a22o_2 _14942_ (.A1(\cpuregs[16][29] ),
    .A2(_11533_),
    .B1(_11451_),
    .B2(_11536_),
    .X(_03340_));
 sky130_fd_sc_hd__a22o_2 _14943_ (.A1(\cpuregs[16][28] ),
    .A2(_11533_),
    .B1(_11452_),
    .B2(_11536_),
    .X(_03339_));
 sky130_fd_sc_hd__a22o_2 _14944_ (.A1(\cpuregs[16][27] ),
    .A2(_11533_),
    .B1(_11453_),
    .B2(_11536_),
    .X(_03338_));
 sky130_fd_sc_hd__a22o_2 _14945_ (.A1(\cpuregs[16][26] ),
    .A2(_11533_),
    .B1(_11454_),
    .B2(_11536_),
    .X(_03337_));
 sky130_fd_sc_hd__buf_1 _14946_ (.A(_11532_),
    .X(_11537_));
 sky130_fd_sc_hd__buf_1 _14947_ (.A(_11535_),
    .X(_11538_));
 sky130_fd_sc_hd__a22o_2 _14948_ (.A1(\cpuregs[16][25] ),
    .A2(_11537_),
    .B1(_11456_),
    .B2(_11538_),
    .X(_03336_));
 sky130_fd_sc_hd__a22o_2 _14949_ (.A1(\cpuregs[16][24] ),
    .A2(_11537_),
    .B1(_11458_),
    .B2(_11538_),
    .X(_03335_));
 sky130_fd_sc_hd__a22o_2 _14950_ (.A1(\cpuregs[16][23] ),
    .A2(_11537_),
    .B1(_11459_),
    .B2(_11538_),
    .X(_03334_));
 sky130_fd_sc_hd__a22o_2 _14951_ (.A1(\cpuregs[16][22] ),
    .A2(_11537_),
    .B1(_11460_),
    .B2(_11538_),
    .X(_03333_));
 sky130_fd_sc_hd__a22o_2 _14952_ (.A1(\cpuregs[16][21] ),
    .A2(_11537_),
    .B1(_11461_),
    .B2(_11538_),
    .X(_03332_));
 sky130_fd_sc_hd__a22o_2 _14953_ (.A1(\cpuregs[16][20] ),
    .A2(_11537_),
    .B1(_11462_),
    .B2(_11538_),
    .X(_03331_));
 sky130_fd_sc_hd__buf_1 _14954_ (.A(_11532_),
    .X(_11539_));
 sky130_fd_sc_hd__buf_1 _14955_ (.A(_11535_),
    .X(_11540_));
 sky130_fd_sc_hd__a22o_2 _14956_ (.A1(\cpuregs[16][19] ),
    .A2(_11539_),
    .B1(_11464_),
    .B2(_11540_),
    .X(_03330_));
 sky130_fd_sc_hd__a22o_2 _14957_ (.A1(\cpuregs[16][18] ),
    .A2(_11539_),
    .B1(_11466_),
    .B2(_11540_),
    .X(_03329_));
 sky130_fd_sc_hd__a22o_2 _14958_ (.A1(\cpuregs[16][17] ),
    .A2(_11539_),
    .B1(_11467_),
    .B2(_11540_),
    .X(_03328_));
 sky130_fd_sc_hd__a22o_2 _14959_ (.A1(\cpuregs[16][16] ),
    .A2(_11539_),
    .B1(_11468_),
    .B2(_11540_),
    .X(_03327_));
 sky130_fd_sc_hd__a22o_2 _14960_ (.A1(\cpuregs[16][15] ),
    .A2(_11539_),
    .B1(_11469_),
    .B2(_11540_),
    .X(_03326_));
 sky130_fd_sc_hd__a22o_2 _14961_ (.A1(\cpuregs[16][14] ),
    .A2(_11539_),
    .B1(_11470_),
    .B2(_11540_),
    .X(_03325_));
 sky130_fd_sc_hd__buf_1 _14962_ (.A(_11532_),
    .X(_11541_));
 sky130_fd_sc_hd__buf_1 _14963_ (.A(_11535_),
    .X(_11542_));
 sky130_fd_sc_hd__a22o_2 _14964_ (.A1(\cpuregs[16][13] ),
    .A2(_11541_),
    .B1(_11472_),
    .B2(_11542_),
    .X(_03324_));
 sky130_fd_sc_hd__a22o_2 _14965_ (.A1(\cpuregs[16][12] ),
    .A2(_11541_),
    .B1(_11474_),
    .B2(_11542_),
    .X(_03323_));
 sky130_fd_sc_hd__a22o_2 _14966_ (.A1(\cpuregs[16][11] ),
    .A2(_11541_),
    .B1(_11475_),
    .B2(_11542_),
    .X(_03322_));
 sky130_fd_sc_hd__a22o_2 _14967_ (.A1(\cpuregs[16][10] ),
    .A2(_11541_),
    .B1(_11476_),
    .B2(_11542_),
    .X(_03321_));
 sky130_fd_sc_hd__a22o_2 _14968_ (.A1(\cpuregs[16][9] ),
    .A2(_11541_),
    .B1(_11477_),
    .B2(_11542_),
    .X(_03320_));
 sky130_fd_sc_hd__a22o_2 _14969_ (.A1(\cpuregs[16][8] ),
    .A2(_11541_),
    .B1(_11478_),
    .B2(_11542_),
    .X(_03319_));
 sky130_fd_sc_hd__buf_1 _14970_ (.A(_11531_),
    .X(_11543_));
 sky130_fd_sc_hd__buf_1 _14971_ (.A(_11534_),
    .X(_11544_));
 sky130_fd_sc_hd__a22o_2 _14972_ (.A1(\cpuregs[16][7] ),
    .A2(_11543_),
    .B1(_11480_),
    .B2(_11544_),
    .X(_03318_));
 sky130_fd_sc_hd__a22o_2 _14973_ (.A1(\cpuregs[16][6] ),
    .A2(_11543_),
    .B1(_11482_),
    .B2(_11544_),
    .X(_03317_));
 sky130_fd_sc_hd__a22o_2 _14974_ (.A1(\cpuregs[16][5] ),
    .A2(_11543_),
    .B1(_11483_),
    .B2(_11544_),
    .X(_03316_));
 sky130_fd_sc_hd__a22o_2 _14975_ (.A1(\cpuregs[16][4] ),
    .A2(_11543_),
    .B1(_11484_),
    .B2(_11544_),
    .X(_03315_));
 sky130_fd_sc_hd__a22o_2 _14976_ (.A1(\cpuregs[16][3] ),
    .A2(_11543_),
    .B1(_11485_),
    .B2(_11544_),
    .X(_03314_));
 sky130_fd_sc_hd__a22o_2 _14977_ (.A1(\cpuregs[16][2] ),
    .A2(_11543_),
    .B1(_11486_),
    .B2(_11544_),
    .X(_03313_));
 sky130_fd_sc_hd__a22o_2 _14978_ (.A1(\cpuregs[16][1] ),
    .A2(_11532_),
    .B1(_11487_),
    .B2(_11535_),
    .X(_03312_));
 sky130_fd_sc_hd__a22o_2 _14979_ (.A1(\cpuregs[16][0] ),
    .A2(_11532_),
    .B1(_11488_),
    .B2(_11535_),
    .X(_03311_));
 sky130_fd_sc_hd__or4_2 _14980_ (.A(_11380_),
    .B(_11310_),
    .C(_11252_),
    .D(_11313_),
    .X(_11545_));
 sky130_fd_sc_hd__buf_1 _14981_ (.A(_11545_),
    .X(_11546_));
 sky130_fd_sc_hd__buf_1 _14982_ (.A(_11546_),
    .X(_11547_));
 sky130_vsdinv _14983_ (.A(_11545_),
    .Y(_11548_));
 sky130_fd_sc_hd__buf_1 _14984_ (.A(_11548_),
    .X(_11549_));
 sky130_fd_sc_hd__buf_1 _14985_ (.A(_11549_),
    .X(_11550_));
 sky130_fd_sc_hd__a22o_2 _14986_ (.A1(\cpuregs[17][31] ),
    .A2(_11547_),
    .B1(_11446_),
    .B2(_11550_),
    .X(_03310_));
 sky130_fd_sc_hd__a22o_2 _14987_ (.A1(\cpuregs[17][30] ),
    .A2(_11547_),
    .B1(_11450_),
    .B2(_11550_),
    .X(_03309_));
 sky130_fd_sc_hd__a22o_2 _14988_ (.A1(\cpuregs[17][29] ),
    .A2(_11547_),
    .B1(_11451_),
    .B2(_11550_),
    .X(_03308_));
 sky130_fd_sc_hd__a22o_2 _14989_ (.A1(\cpuregs[17][28] ),
    .A2(_11547_),
    .B1(_11452_),
    .B2(_11550_),
    .X(_03307_));
 sky130_fd_sc_hd__a22o_2 _14990_ (.A1(\cpuregs[17][27] ),
    .A2(_11547_),
    .B1(_11453_),
    .B2(_11550_),
    .X(_03306_));
 sky130_fd_sc_hd__a22o_2 _14991_ (.A1(\cpuregs[17][26] ),
    .A2(_11547_),
    .B1(_11454_),
    .B2(_11550_),
    .X(_03305_));
 sky130_fd_sc_hd__buf_1 _14992_ (.A(_11546_),
    .X(_11551_));
 sky130_fd_sc_hd__buf_1 _14993_ (.A(_11549_),
    .X(_11552_));
 sky130_fd_sc_hd__a22o_2 _14994_ (.A1(\cpuregs[17][25] ),
    .A2(_11551_),
    .B1(_11456_),
    .B2(_11552_),
    .X(_03304_));
 sky130_fd_sc_hd__a22o_2 _14995_ (.A1(\cpuregs[17][24] ),
    .A2(_11551_),
    .B1(_11458_),
    .B2(_11552_),
    .X(_03303_));
 sky130_fd_sc_hd__a22o_2 _14996_ (.A1(\cpuregs[17][23] ),
    .A2(_11551_),
    .B1(_11459_),
    .B2(_11552_),
    .X(_03302_));
 sky130_fd_sc_hd__a22o_2 _14997_ (.A1(\cpuregs[17][22] ),
    .A2(_11551_),
    .B1(_11460_),
    .B2(_11552_),
    .X(_03301_));
 sky130_fd_sc_hd__a22o_2 _14998_ (.A1(\cpuregs[17][21] ),
    .A2(_11551_),
    .B1(_11461_),
    .B2(_11552_),
    .X(_03300_));
 sky130_fd_sc_hd__a22o_2 _14999_ (.A1(\cpuregs[17][20] ),
    .A2(_11551_),
    .B1(_11462_),
    .B2(_11552_),
    .X(_03299_));
 sky130_fd_sc_hd__buf_1 _15000_ (.A(_11546_),
    .X(_11553_));
 sky130_fd_sc_hd__buf_1 _15001_ (.A(_11549_),
    .X(_11554_));
 sky130_fd_sc_hd__a22o_2 _15002_ (.A1(\cpuregs[17][19] ),
    .A2(_11553_),
    .B1(_11464_),
    .B2(_11554_),
    .X(_03298_));
 sky130_fd_sc_hd__a22o_2 _15003_ (.A1(\cpuregs[17][18] ),
    .A2(_11553_),
    .B1(_11466_),
    .B2(_11554_),
    .X(_03297_));
 sky130_fd_sc_hd__a22o_2 _15004_ (.A1(\cpuregs[17][17] ),
    .A2(_11553_),
    .B1(_11467_),
    .B2(_11554_),
    .X(_03296_));
 sky130_fd_sc_hd__a22o_2 _15005_ (.A1(\cpuregs[17][16] ),
    .A2(_11553_),
    .B1(_11468_),
    .B2(_11554_),
    .X(_03295_));
 sky130_fd_sc_hd__a22o_2 _15006_ (.A1(\cpuregs[17][15] ),
    .A2(_11553_),
    .B1(_11469_),
    .B2(_11554_),
    .X(_03294_));
 sky130_fd_sc_hd__a22o_2 _15007_ (.A1(\cpuregs[17][14] ),
    .A2(_11553_),
    .B1(_11470_),
    .B2(_11554_),
    .X(_03293_));
 sky130_fd_sc_hd__buf_1 _15008_ (.A(_11546_),
    .X(_11555_));
 sky130_fd_sc_hd__buf_1 _15009_ (.A(_11549_),
    .X(_11556_));
 sky130_fd_sc_hd__a22o_2 _15010_ (.A1(\cpuregs[17][13] ),
    .A2(_11555_),
    .B1(_11472_),
    .B2(_11556_),
    .X(_03292_));
 sky130_fd_sc_hd__a22o_2 _15011_ (.A1(\cpuregs[17][12] ),
    .A2(_11555_),
    .B1(_11474_),
    .B2(_11556_),
    .X(_03291_));
 sky130_fd_sc_hd__a22o_2 _15012_ (.A1(\cpuregs[17][11] ),
    .A2(_11555_),
    .B1(_11475_),
    .B2(_11556_),
    .X(_03290_));
 sky130_fd_sc_hd__a22o_2 _15013_ (.A1(\cpuregs[17][10] ),
    .A2(_11555_),
    .B1(_11476_),
    .B2(_11556_),
    .X(_03289_));
 sky130_fd_sc_hd__a22o_2 _15014_ (.A1(\cpuregs[17][9] ),
    .A2(_11555_),
    .B1(_11477_),
    .B2(_11556_),
    .X(_03288_));
 sky130_fd_sc_hd__a22o_2 _15015_ (.A1(\cpuregs[17][8] ),
    .A2(_11555_),
    .B1(_11478_),
    .B2(_11556_),
    .X(_03287_));
 sky130_fd_sc_hd__buf_1 _15016_ (.A(_11545_),
    .X(_11557_));
 sky130_fd_sc_hd__buf_1 _15017_ (.A(_11548_),
    .X(_11558_));
 sky130_fd_sc_hd__a22o_2 _15018_ (.A1(\cpuregs[17][7] ),
    .A2(_11557_),
    .B1(_11480_),
    .B2(_11558_),
    .X(_03286_));
 sky130_fd_sc_hd__a22o_2 _15019_ (.A1(\cpuregs[17][6] ),
    .A2(_11557_),
    .B1(_11482_),
    .B2(_11558_),
    .X(_03285_));
 sky130_fd_sc_hd__a22o_2 _15020_ (.A1(\cpuregs[17][5] ),
    .A2(_11557_),
    .B1(_11483_),
    .B2(_11558_),
    .X(_03284_));
 sky130_fd_sc_hd__a22o_2 _15021_ (.A1(\cpuregs[17][4] ),
    .A2(_11557_),
    .B1(_11484_),
    .B2(_11558_),
    .X(_03283_));
 sky130_fd_sc_hd__a22o_2 _15022_ (.A1(\cpuregs[17][3] ),
    .A2(_11557_),
    .B1(_11485_),
    .B2(_11558_),
    .X(_03282_));
 sky130_fd_sc_hd__a22o_2 _15023_ (.A1(\cpuregs[17][2] ),
    .A2(_11557_),
    .B1(_11486_),
    .B2(_11558_),
    .X(_03281_));
 sky130_fd_sc_hd__a22o_2 _15024_ (.A1(\cpuregs[17][1] ),
    .A2(_11546_),
    .B1(_11487_),
    .B2(_11549_),
    .X(_03280_));
 sky130_fd_sc_hd__a22o_2 _15025_ (.A1(\cpuregs[17][0] ),
    .A2(_11546_),
    .B1(_11488_),
    .B2(_11549_),
    .X(_03279_));
 sky130_fd_sc_hd__buf_1 _15026_ (.A(\pcpi_mul.rs2[31] ),
    .X(_11559_));
 sky130_fd_sc_hd__buf_1 _15027_ (.A(_11559_),
    .X(_11560_));
 sky130_fd_sc_hd__buf_1 _15028_ (.A(_11560_),
    .X(_11561_));
 sky130_fd_sc_hd__buf_1 _15029_ (.A(_11561_),
    .X(_11562_));
 sky130_fd_sc_hd__buf_1 _15030_ (.A(_11562_),
    .X(_11563_));
 sky130_fd_sc_hd__buf_1 _15031_ (.A(_10578_),
    .X(_11564_));
 sky130_fd_sc_hd__buf_1 _15032_ (.A(_11564_),
    .X(_11565_));
 sky130_fd_sc_hd__a22o_2 _15033_ (.A1(pcpi_rs2[31]),
    .A2(_10592_),
    .B1(_11563_),
    .B2(_11565_),
    .X(_03278_));
 sky130_fd_sc_hd__a22o_2 _15034_ (.A1(\pcpi_mul.rs2[30] ),
    .A2(_11565_),
    .B1(pcpi_rs2[30]),
    .B2(_03728_),
    .X(_03277_));
 sky130_fd_sc_hd__buf_1 _15035_ (.A(\pcpi_mul.rs2[29] ),
    .X(_11566_));
 sky130_fd_sc_hd__buf_1 _15036_ (.A(_11566_),
    .X(_11567_));
 sky130_fd_sc_hd__buf_1 _15037_ (.A(_11567_),
    .X(_11568_));
 sky130_fd_sc_hd__buf_1 _15038_ (.A(_11568_),
    .X(_11569_));
 sky130_fd_sc_hd__a22o_2 _15039_ (.A1(_11569_),
    .A2(_11565_),
    .B1(_11334_),
    .B2(_03728_),
    .X(_03276_));
 sky130_fd_sc_hd__buf_1 _15040_ (.A(\pcpi_mul.rs2[28] ),
    .X(_11570_));
 sky130_fd_sc_hd__buf_1 _15041_ (.A(_11570_),
    .X(_11571_));
 sky130_fd_sc_hd__buf_1 _15042_ (.A(_11571_),
    .X(_11572_));
 sky130_fd_sc_hd__buf_1 _15043_ (.A(_11572_),
    .X(_11573_));
 sky130_fd_sc_hd__a22o_2 _15044_ (.A1(_11573_),
    .A2(_11565_),
    .B1(pcpi_rs2[28]),
    .B2(_03728_),
    .X(_03275_));
 sky130_fd_sc_hd__a22o_2 _15045_ (.A1(\pcpi_mul.rs2[27] ),
    .A2(_11565_),
    .B1(_11335_),
    .B2(_03728_),
    .X(_03274_));
 sky130_fd_sc_hd__buf_1 _15046_ (.A(\pcpi_mul.rs2[26] ),
    .X(_11574_));
 sky130_fd_sc_hd__buf_1 _15047_ (.A(_11574_),
    .X(_11575_));
 sky130_fd_sc_hd__buf_1 _15048_ (.A(_11575_),
    .X(_11576_));
 sky130_fd_sc_hd__buf_1 _15049_ (.A(_11576_),
    .X(_11577_));
 sky130_fd_sc_hd__buf_1 _15050_ (.A(_11564_),
    .X(_11578_));
 sky130_fd_sc_hd__a22o_2 _15051_ (.A1(_11577_),
    .A2(_11578_),
    .B1(pcpi_rs2[26]),
    .B2(_03728_),
    .X(_03273_));
 sky130_fd_sc_hd__buf_1 _15052_ (.A(\pcpi_mul.rs2[25] ),
    .X(_11579_));
 sky130_fd_sc_hd__buf_1 _15053_ (.A(_11579_),
    .X(_11580_));
 sky130_fd_sc_hd__buf_1 _15054_ (.A(_11580_),
    .X(_11581_));
 sky130_fd_sc_hd__buf_1 _15055_ (.A(_11581_),
    .X(_11582_));
 sky130_fd_sc_hd__buf_1 _15056_ (.A(_10601_),
    .X(_11583_));
 sky130_fd_sc_hd__a22o_2 _15057_ (.A1(_11582_),
    .A2(_11578_),
    .B1(_11337_),
    .B2(_11583_),
    .X(_03272_));
 sky130_fd_sc_hd__a22o_2 _15058_ (.A1(\pcpi_mul.rs2[24] ),
    .A2(_11578_),
    .B1(pcpi_rs2[24]),
    .B2(_11583_),
    .X(_03271_));
 sky130_fd_sc_hd__buf_1 _15059_ (.A(\pcpi_mul.rs2[23] ),
    .X(_11584_));
 sky130_fd_sc_hd__buf_1 _15060_ (.A(_11584_),
    .X(_11585_));
 sky130_fd_sc_hd__buf_1 _15061_ (.A(_11585_),
    .X(_11586_));
 sky130_fd_sc_hd__buf_1 _15062_ (.A(_11586_),
    .X(_11587_));
 sky130_fd_sc_hd__a22o_2 _15063_ (.A1(_11587_),
    .A2(_11578_),
    .B1(_11339_),
    .B2(_11583_),
    .X(_03270_));
 sky130_fd_sc_hd__buf_1 _15064_ (.A(\pcpi_mul.rs2[22] ),
    .X(_11588_));
 sky130_fd_sc_hd__buf_1 _15065_ (.A(_11588_),
    .X(_11589_));
 sky130_fd_sc_hd__buf_1 _15066_ (.A(_11589_),
    .X(_11590_));
 sky130_fd_sc_hd__buf_1 _15067_ (.A(_11590_),
    .X(_11591_));
 sky130_fd_sc_hd__a22o_2 _15068_ (.A1(_11591_),
    .A2(_11578_),
    .B1(pcpi_rs2[22]),
    .B2(_11583_),
    .X(_03269_));
 sky130_fd_sc_hd__a22o_2 _15069_ (.A1(\pcpi_mul.rs2[21] ),
    .A2(_11578_),
    .B1(_11340_),
    .B2(_11583_),
    .X(_03268_));
 sky130_fd_sc_hd__buf_1 _15070_ (.A(\pcpi_mul.rs2[20] ),
    .X(_11592_));
 sky130_fd_sc_hd__buf_1 _15071_ (.A(_11592_),
    .X(_11593_));
 sky130_fd_sc_hd__buf_1 _15072_ (.A(_11593_),
    .X(_11594_));
 sky130_fd_sc_hd__buf_1 _15073_ (.A(_10578_),
    .X(_11595_));
 sky130_fd_sc_hd__buf_1 _15074_ (.A(_11595_),
    .X(_11596_));
 sky130_fd_sc_hd__a22o_2 _15075_ (.A1(_11594_),
    .A2(_11596_),
    .B1(pcpi_rs2[20]),
    .B2(_11583_),
    .X(_03267_));
 sky130_fd_sc_hd__buf_1 _15076_ (.A(\pcpi_mul.rs2[19] ),
    .X(_11597_));
 sky130_fd_sc_hd__buf_1 _15077_ (.A(_11597_),
    .X(_11598_));
 sky130_fd_sc_hd__buf_1 _15078_ (.A(_11598_),
    .X(_11599_));
 sky130_fd_sc_hd__buf_1 _15079_ (.A(_10601_),
    .X(_11600_));
 sky130_fd_sc_hd__a22o_2 _15080_ (.A1(_11599_),
    .A2(_11596_),
    .B1(_11342_),
    .B2(_11600_),
    .X(_03266_));
 sky130_fd_sc_hd__a22o_2 _15081_ (.A1(\pcpi_mul.rs2[18] ),
    .A2(_11596_),
    .B1(pcpi_rs2[18]),
    .B2(_11600_),
    .X(_03265_));
 sky130_fd_sc_hd__buf_1 _15082_ (.A(\pcpi_mul.rs2[17] ),
    .X(_11601_));
 sky130_fd_sc_hd__buf_1 _15083_ (.A(_11601_),
    .X(_11602_));
 sky130_fd_sc_hd__buf_1 _15084_ (.A(_11602_),
    .X(_11603_));
 sky130_fd_sc_hd__a22o_2 _15085_ (.A1(_11603_),
    .A2(_11596_),
    .B1(_11344_),
    .B2(_11600_),
    .X(_03264_));
 sky130_fd_sc_hd__buf_1 _15086_ (.A(\pcpi_mul.rs2[16] ),
    .X(_11604_));
 sky130_fd_sc_hd__buf_1 _15087_ (.A(_11604_),
    .X(_11605_));
 sky130_fd_sc_hd__buf_1 _15088_ (.A(_11605_),
    .X(_11606_));
 sky130_fd_sc_hd__a22o_2 _15089_ (.A1(_11606_),
    .A2(_11596_),
    .B1(pcpi_rs2[16]),
    .B2(_11600_),
    .X(_03263_));
 sky130_fd_sc_hd__a22o_2 _15090_ (.A1(\pcpi_mul.rs2[15] ),
    .A2(_11596_),
    .B1(_11345_),
    .B2(_11600_),
    .X(_03262_));
 sky130_fd_sc_hd__buf_1 _15091_ (.A(\pcpi_mul.rs2[14] ),
    .X(_11607_));
 sky130_fd_sc_hd__buf_1 _15092_ (.A(_11607_),
    .X(_11608_));
 sky130_fd_sc_hd__buf_1 _15093_ (.A(_11595_),
    .X(_11609_));
 sky130_fd_sc_hd__a22o_2 _15094_ (.A1(_11608_),
    .A2(_11609_),
    .B1(_11346_),
    .B2(_11600_),
    .X(_03261_));
 sky130_fd_sc_hd__buf_1 _15095_ (.A(\pcpi_mul.rs2[13] ),
    .X(_11610_));
 sky130_fd_sc_hd__buf_1 _15096_ (.A(_11610_),
    .X(_11611_));
 sky130_fd_sc_hd__buf_1 _15097_ (.A(_10601_),
    .X(_11612_));
 sky130_fd_sc_hd__a22o_2 _15098_ (.A1(_11611_),
    .A2(_11609_),
    .B1(_11348_),
    .B2(_11612_),
    .X(_03260_));
 sky130_fd_sc_hd__a22o_2 _15099_ (.A1(\pcpi_mul.rs2[12] ),
    .A2(_11609_),
    .B1(_11350_),
    .B2(_11612_),
    .X(_03259_));
 sky130_fd_sc_hd__buf_1 _15100_ (.A(\pcpi_mul.rs2[11] ),
    .X(_11613_));
 sky130_fd_sc_hd__buf_1 _15101_ (.A(_11613_),
    .X(_11614_));
 sky130_fd_sc_hd__a22o_2 _15102_ (.A1(_11614_),
    .A2(_11609_),
    .B1(_11351_),
    .B2(_11612_),
    .X(_03258_));
 sky130_fd_sc_hd__buf_1 _15103_ (.A(\pcpi_mul.rs2[10] ),
    .X(_11615_));
 sky130_fd_sc_hd__buf_1 _15104_ (.A(_11615_),
    .X(_11616_));
 sky130_fd_sc_hd__buf_1 _15105_ (.A(_11616_),
    .X(_11617_));
 sky130_fd_sc_hd__a22o_2 _15106_ (.A1(_11617_),
    .A2(_11609_),
    .B1(_11352_),
    .B2(_11612_),
    .X(_03257_));
 sky130_fd_sc_hd__a22o_2 _15107_ (.A1(\pcpi_mul.rs2[9] ),
    .A2(_11609_),
    .B1(_11353_),
    .B2(_11612_),
    .X(_03256_));
 sky130_fd_sc_hd__buf_1 _15108_ (.A(\pcpi_mul.rs2[8] ),
    .X(_11618_));
 sky130_fd_sc_hd__buf_1 _15109_ (.A(_11618_),
    .X(_11619_));
 sky130_fd_sc_hd__buf_1 _15110_ (.A(_11619_),
    .X(_11620_));
 sky130_fd_sc_hd__buf_1 _15111_ (.A(_11595_),
    .X(_11621_));
 sky130_fd_sc_hd__a22o_2 _15112_ (.A1(_11620_),
    .A2(_11621_),
    .B1(_11354_),
    .B2(_11612_),
    .X(_03255_));
 sky130_fd_sc_hd__buf_1 _15113_ (.A(\pcpi_mul.rs2[7] ),
    .X(_11622_));
 sky130_fd_sc_hd__buf_1 _15114_ (.A(_11622_),
    .X(_11623_));
 sky130_fd_sc_hd__buf_1 _15115_ (.A(_11623_),
    .X(_11624_));
 sky130_fd_sc_hd__buf_1 _15116_ (.A(_10601_),
    .X(_11625_));
 sky130_fd_sc_hd__a22o_2 _15117_ (.A1(_11624_),
    .A2(_11621_),
    .B1(_11356_),
    .B2(_11625_),
    .X(_03254_));
 sky130_fd_sc_hd__a22o_2 _15118_ (.A1(\pcpi_mul.rs2[6] ),
    .A2(_11621_),
    .B1(_11358_),
    .B2(_11625_),
    .X(_03253_));
 sky130_fd_sc_hd__buf_1 _15119_ (.A(\pcpi_mul.rs2[5] ),
    .X(_11626_));
 sky130_fd_sc_hd__buf_1 _15120_ (.A(_11626_),
    .X(_11627_));
 sky130_fd_sc_hd__buf_1 _15121_ (.A(_11627_),
    .X(_11628_));
 sky130_fd_sc_hd__buf_1 _15122_ (.A(_11628_),
    .X(_11629_));
 sky130_fd_sc_hd__a22o_2 _15123_ (.A1(_11629_),
    .A2(_11621_),
    .B1(_11359_),
    .B2(_11625_),
    .X(_03252_));
 sky130_fd_sc_hd__buf_1 _15124_ (.A(\pcpi_mul.rs2[4] ),
    .X(_11630_));
 sky130_fd_sc_hd__buf_1 _15125_ (.A(_11630_),
    .X(_11631_));
 sky130_fd_sc_hd__buf_1 _15126_ (.A(_11631_),
    .X(_11632_));
 sky130_fd_sc_hd__buf_1 _15127_ (.A(_11632_),
    .X(_11633_));
 sky130_fd_sc_hd__a22o_2 _15128_ (.A1(_11633_),
    .A2(_11621_),
    .B1(_11360_),
    .B2(_11625_),
    .X(_03251_));
 sky130_fd_sc_hd__a22o_2 _15129_ (.A1(\pcpi_mul.rs2[3] ),
    .A2(_11621_),
    .B1(_11361_),
    .B2(_11625_),
    .X(_03250_));
 sky130_fd_sc_hd__buf_1 _15130_ (.A(\pcpi_mul.rs2[2] ),
    .X(_11634_));
 sky130_fd_sc_hd__buf_1 _15131_ (.A(_11634_),
    .X(_11635_));
 sky130_fd_sc_hd__buf_1 _15132_ (.A(_11635_),
    .X(_11636_));
 sky130_fd_sc_hd__buf_1 _15133_ (.A(_11636_),
    .X(_11637_));
 sky130_fd_sc_hd__buf_1 _15134_ (.A(_11637_),
    .X(_11638_));
 sky130_fd_sc_hd__buf_1 _15135_ (.A(_11595_),
    .X(_11639_));
 sky130_fd_sc_hd__a22o_2 _15136_ (.A1(_11638_),
    .A2(_11639_),
    .B1(_11362_),
    .B2(_11625_),
    .X(_03249_));
 sky130_fd_sc_hd__buf_1 _15137_ (.A(\pcpi_mul.rs2[1] ),
    .X(_11640_));
 sky130_fd_sc_hd__buf_1 _15138_ (.A(_11640_),
    .X(_11641_));
 sky130_fd_sc_hd__buf_1 _15139_ (.A(_11641_),
    .X(_11642_));
 sky130_fd_sc_hd__buf_1 _15140_ (.A(_11642_),
    .X(_11643_));
 sky130_fd_sc_hd__buf_1 _15141_ (.A(_11643_),
    .X(_11644_));
 sky130_fd_sc_hd__buf_1 _15142_ (.A(_10591_),
    .X(_11645_));
 sky130_fd_sc_hd__a22o_2 _15143_ (.A1(_11644_),
    .A2(_11639_),
    .B1(_11363_),
    .B2(_11645_),
    .X(_03248_));
 sky130_fd_sc_hd__a22o_2 _15144_ (.A1(\pcpi_mul.rs2[0] ),
    .A2(_11639_),
    .B1(_11364_),
    .B2(_11645_),
    .X(_03247_));
 sky130_fd_sc_hd__a22o_2 _15145_ (.A1(mem_wstrb[3]),
    .A2(_10478_),
    .B1(_02541_),
    .B2(_10480_),
    .X(_03246_));
 sky130_fd_sc_hd__a22o_2 _15146_ (.A1(mem_wstrb[2]),
    .A2(_10478_),
    .B1(_02540_),
    .B2(_10480_),
    .X(_03245_));
 sky130_fd_sc_hd__a22o_2 _15147_ (.A1(mem_wstrb[1]),
    .A2(_10478_),
    .B1(_02539_),
    .B2(_10480_),
    .X(_03244_));
 sky130_fd_sc_hd__a22o_2 _15148_ (.A1(mem_wstrb[0]),
    .A2(_10478_),
    .B1(_02538_),
    .B2(_10480_),
    .X(_03243_));
 sky130_vsdinv _15149_ (.A(_10714_),
    .Y(_11646_));
 sky130_fd_sc_hd__or4_2 _15150_ (.A(_00327_),
    .B(_10499_),
    .C(_00330_),
    .D(_10491_),
    .X(_11647_));
 sky130_fd_sc_hd__o32a_2 _15151_ (.A1(_10713_),
    .A2(_11646_),
    .A3(_11647_),
    .B1(_10730_),
    .B2(_10506_),
    .X(_11648_));
 sky130_vsdinv _15152_ (.A(_11648_),
    .Y(_03242_));
 sky130_fd_sc_hd__o32a_2 _15153_ (.A1(_00329_),
    .A2(_11646_),
    .A3(_11647_),
    .B1(_10769_),
    .B2(_10493_),
    .X(_11649_));
 sky130_vsdinv _15154_ (.A(_11649_),
    .Y(_03241_));
 sky130_fd_sc_hd__or2_2 _15155_ (.A(_11313_),
    .B(_11428_),
    .X(_11650_));
 sky130_fd_sc_hd__buf_1 _15156_ (.A(_11650_),
    .X(_11651_));
 sky130_fd_sc_hd__buf_1 _15157_ (.A(_11651_),
    .X(_11652_));
 sky130_fd_sc_hd__buf_1 _15158_ (.A(\cpuregs_wrdata[31] ),
    .X(_11653_));
 sky130_vsdinv _15159_ (.A(_11650_),
    .Y(_11654_));
 sky130_fd_sc_hd__buf_1 _15160_ (.A(_11654_),
    .X(_11655_));
 sky130_fd_sc_hd__buf_1 _15161_ (.A(_11655_),
    .X(_11656_));
 sky130_fd_sc_hd__a22o_2 _15162_ (.A1(\cpuregs[13][31] ),
    .A2(_11652_),
    .B1(_11653_),
    .B2(_11656_),
    .X(_03240_));
 sky130_fd_sc_hd__buf_1 _15163_ (.A(\cpuregs_wrdata[30] ),
    .X(_11657_));
 sky130_fd_sc_hd__a22o_2 _15164_ (.A1(\cpuregs[13][30] ),
    .A2(_11652_),
    .B1(_11657_),
    .B2(_11656_),
    .X(_03239_));
 sky130_fd_sc_hd__buf_1 _15165_ (.A(\cpuregs_wrdata[29] ),
    .X(_11658_));
 sky130_fd_sc_hd__a22o_2 _15166_ (.A1(\cpuregs[13][29] ),
    .A2(_11652_),
    .B1(_11658_),
    .B2(_11656_),
    .X(_03238_));
 sky130_fd_sc_hd__buf_1 _15167_ (.A(\cpuregs_wrdata[28] ),
    .X(_11659_));
 sky130_fd_sc_hd__a22o_2 _15168_ (.A1(\cpuregs[13][28] ),
    .A2(_11652_),
    .B1(_11659_),
    .B2(_11656_),
    .X(_03237_));
 sky130_fd_sc_hd__buf_1 _15169_ (.A(\cpuregs_wrdata[27] ),
    .X(_11660_));
 sky130_fd_sc_hd__a22o_2 _15170_ (.A1(\cpuregs[13][27] ),
    .A2(_11652_),
    .B1(_11660_),
    .B2(_11656_),
    .X(_03236_));
 sky130_fd_sc_hd__buf_1 _15171_ (.A(\cpuregs_wrdata[26] ),
    .X(_11661_));
 sky130_fd_sc_hd__a22o_2 _15172_ (.A1(\cpuregs[13][26] ),
    .A2(_11652_),
    .B1(_11661_),
    .B2(_11656_),
    .X(_03235_));
 sky130_fd_sc_hd__buf_1 _15173_ (.A(_11651_),
    .X(_11662_));
 sky130_fd_sc_hd__buf_1 _15174_ (.A(\cpuregs_wrdata[25] ),
    .X(_11663_));
 sky130_fd_sc_hd__buf_1 _15175_ (.A(_11655_),
    .X(_11664_));
 sky130_fd_sc_hd__a22o_2 _15176_ (.A1(\cpuregs[13][25] ),
    .A2(_11662_),
    .B1(_11663_),
    .B2(_11664_),
    .X(_03234_));
 sky130_fd_sc_hd__buf_1 _15177_ (.A(\cpuregs_wrdata[24] ),
    .X(_11665_));
 sky130_fd_sc_hd__a22o_2 _15178_ (.A1(\cpuregs[13][24] ),
    .A2(_11662_),
    .B1(_11665_),
    .B2(_11664_),
    .X(_03233_));
 sky130_fd_sc_hd__buf_1 _15179_ (.A(\cpuregs_wrdata[23] ),
    .X(_11666_));
 sky130_fd_sc_hd__a22o_2 _15180_ (.A1(\cpuregs[13][23] ),
    .A2(_11662_),
    .B1(_11666_),
    .B2(_11664_),
    .X(_03232_));
 sky130_fd_sc_hd__buf_1 _15181_ (.A(\cpuregs_wrdata[22] ),
    .X(_11667_));
 sky130_fd_sc_hd__a22o_2 _15182_ (.A1(\cpuregs[13][22] ),
    .A2(_11662_),
    .B1(_11667_),
    .B2(_11664_),
    .X(_03231_));
 sky130_fd_sc_hd__buf_1 _15183_ (.A(\cpuregs_wrdata[21] ),
    .X(_11668_));
 sky130_fd_sc_hd__a22o_2 _15184_ (.A1(\cpuregs[13][21] ),
    .A2(_11662_),
    .B1(_11668_),
    .B2(_11664_),
    .X(_03230_));
 sky130_fd_sc_hd__buf_1 _15185_ (.A(\cpuregs_wrdata[20] ),
    .X(_11669_));
 sky130_fd_sc_hd__a22o_2 _15186_ (.A1(\cpuregs[13][20] ),
    .A2(_11662_),
    .B1(_11669_),
    .B2(_11664_),
    .X(_03229_));
 sky130_fd_sc_hd__buf_1 _15187_ (.A(_11651_),
    .X(_11670_));
 sky130_fd_sc_hd__buf_1 _15188_ (.A(\cpuregs_wrdata[19] ),
    .X(_11671_));
 sky130_fd_sc_hd__buf_1 _15189_ (.A(_11655_),
    .X(_11672_));
 sky130_fd_sc_hd__a22o_2 _15190_ (.A1(\cpuregs[13][19] ),
    .A2(_11670_),
    .B1(_11671_),
    .B2(_11672_),
    .X(_03228_));
 sky130_fd_sc_hd__buf_1 _15191_ (.A(\cpuregs_wrdata[18] ),
    .X(_11673_));
 sky130_fd_sc_hd__a22o_2 _15192_ (.A1(\cpuregs[13][18] ),
    .A2(_11670_),
    .B1(_11673_),
    .B2(_11672_),
    .X(_03227_));
 sky130_fd_sc_hd__buf_1 _15193_ (.A(\cpuregs_wrdata[17] ),
    .X(_11674_));
 sky130_fd_sc_hd__a22o_2 _15194_ (.A1(\cpuregs[13][17] ),
    .A2(_11670_),
    .B1(_11674_),
    .B2(_11672_),
    .X(_03226_));
 sky130_fd_sc_hd__buf_1 _15195_ (.A(\cpuregs_wrdata[16] ),
    .X(_11675_));
 sky130_fd_sc_hd__a22o_2 _15196_ (.A1(\cpuregs[13][16] ),
    .A2(_11670_),
    .B1(_11675_),
    .B2(_11672_),
    .X(_03225_));
 sky130_fd_sc_hd__buf_1 _15197_ (.A(\cpuregs_wrdata[15] ),
    .X(_11676_));
 sky130_fd_sc_hd__a22o_2 _15198_ (.A1(\cpuregs[13][15] ),
    .A2(_11670_),
    .B1(_11676_),
    .B2(_11672_),
    .X(_03224_));
 sky130_fd_sc_hd__buf_1 _15199_ (.A(\cpuregs_wrdata[14] ),
    .X(_11677_));
 sky130_fd_sc_hd__a22o_2 _15200_ (.A1(\cpuregs[13][14] ),
    .A2(_11670_),
    .B1(_11677_),
    .B2(_11672_),
    .X(_03223_));
 sky130_fd_sc_hd__buf_1 _15201_ (.A(_11651_),
    .X(_11678_));
 sky130_fd_sc_hd__buf_1 _15202_ (.A(\cpuregs_wrdata[13] ),
    .X(_11679_));
 sky130_fd_sc_hd__buf_1 _15203_ (.A(_11655_),
    .X(_11680_));
 sky130_fd_sc_hd__a22o_2 _15204_ (.A1(\cpuregs[13][13] ),
    .A2(_11678_),
    .B1(_11679_),
    .B2(_11680_),
    .X(_03222_));
 sky130_fd_sc_hd__buf_1 _15205_ (.A(\cpuregs_wrdata[12] ),
    .X(_11681_));
 sky130_fd_sc_hd__a22o_2 _15206_ (.A1(\cpuregs[13][12] ),
    .A2(_11678_),
    .B1(_11681_),
    .B2(_11680_),
    .X(_03221_));
 sky130_fd_sc_hd__buf_1 _15207_ (.A(\cpuregs_wrdata[11] ),
    .X(_11682_));
 sky130_fd_sc_hd__a22o_2 _15208_ (.A1(\cpuregs[13][11] ),
    .A2(_11678_),
    .B1(_11682_),
    .B2(_11680_),
    .X(_03220_));
 sky130_fd_sc_hd__buf_1 _15209_ (.A(\cpuregs_wrdata[10] ),
    .X(_11683_));
 sky130_fd_sc_hd__a22o_2 _15210_ (.A1(\cpuregs[13][10] ),
    .A2(_11678_),
    .B1(_11683_),
    .B2(_11680_),
    .X(_03219_));
 sky130_fd_sc_hd__buf_1 _15211_ (.A(\cpuregs_wrdata[9] ),
    .X(_11684_));
 sky130_fd_sc_hd__a22o_2 _15212_ (.A1(\cpuregs[13][9] ),
    .A2(_11678_),
    .B1(_11684_),
    .B2(_11680_),
    .X(_03218_));
 sky130_fd_sc_hd__buf_1 _15213_ (.A(\cpuregs_wrdata[8] ),
    .X(_11685_));
 sky130_fd_sc_hd__a22o_2 _15214_ (.A1(\cpuregs[13][8] ),
    .A2(_11678_),
    .B1(_11685_),
    .B2(_11680_),
    .X(_03217_));
 sky130_fd_sc_hd__buf_1 _15215_ (.A(_11650_),
    .X(_11686_));
 sky130_fd_sc_hd__buf_1 _15216_ (.A(\cpuregs_wrdata[7] ),
    .X(_11687_));
 sky130_fd_sc_hd__buf_1 _15217_ (.A(_11654_),
    .X(_11688_));
 sky130_fd_sc_hd__a22o_2 _15218_ (.A1(\cpuregs[13][7] ),
    .A2(_11686_),
    .B1(_11687_),
    .B2(_11688_),
    .X(_03216_));
 sky130_fd_sc_hd__buf_1 _15219_ (.A(\cpuregs_wrdata[6] ),
    .X(_11689_));
 sky130_fd_sc_hd__a22o_2 _15220_ (.A1(\cpuregs[13][6] ),
    .A2(_11686_),
    .B1(_11689_),
    .B2(_11688_),
    .X(_03215_));
 sky130_fd_sc_hd__buf_1 _15221_ (.A(\cpuregs_wrdata[5] ),
    .X(_11690_));
 sky130_fd_sc_hd__a22o_2 _15222_ (.A1(\cpuregs[13][5] ),
    .A2(_11686_),
    .B1(_11690_),
    .B2(_11688_),
    .X(_03214_));
 sky130_fd_sc_hd__buf_1 _15223_ (.A(\cpuregs_wrdata[4] ),
    .X(_11691_));
 sky130_fd_sc_hd__a22o_2 _15224_ (.A1(\cpuregs[13][4] ),
    .A2(_11686_),
    .B1(_11691_),
    .B2(_11688_),
    .X(_03213_));
 sky130_fd_sc_hd__buf_1 _15225_ (.A(\cpuregs_wrdata[3] ),
    .X(_11692_));
 sky130_fd_sc_hd__a22o_2 _15226_ (.A1(\cpuregs[13][3] ),
    .A2(_11686_),
    .B1(_11692_),
    .B2(_11688_),
    .X(_03212_));
 sky130_fd_sc_hd__buf_1 _15227_ (.A(\cpuregs_wrdata[2] ),
    .X(_11693_));
 sky130_fd_sc_hd__a22o_2 _15228_ (.A1(\cpuregs[13][2] ),
    .A2(_11686_),
    .B1(_11693_),
    .B2(_11688_),
    .X(_03211_));
 sky130_fd_sc_hd__buf_1 _15229_ (.A(\cpuregs_wrdata[1] ),
    .X(_11694_));
 sky130_fd_sc_hd__a22o_2 _15230_ (.A1(\cpuregs[13][1] ),
    .A2(_11651_),
    .B1(_11694_),
    .B2(_11655_),
    .X(_03210_));
 sky130_fd_sc_hd__buf_1 _15231_ (.A(\cpuregs_wrdata[0] ),
    .X(_11695_));
 sky130_fd_sc_hd__a22o_2 _15232_ (.A1(\cpuregs[13][0] ),
    .A2(_11651_),
    .B1(_11695_),
    .B2(_11655_),
    .X(_03209_));
 sky130_fd_sc_hd__o32a_2 _15233_ (.A1(_10713_),
    .A2(_10714_),
    .A3(_11647_),
    .B1(_10666_),
    .B2(_10493_),
    .X(_11696_));
 sky130_vsdinv _15234_ (.A(_11696_),
    .Y(_03208_));
 sky130_fd_sc_hd__a31oi_2 _15235_ (.A1(_00335_),
    .A2(_10756_),
    .A3(_10758_),
    .B1(_10769_),
    .Y(_11697_));
 sky130_fd_sc_hd__buf_1 _15236_ (.A(_10748_),
    .X(_11698_));
 sky130_fd_sc_hd__buf_1 _15237_ (.A(_11698_),
    .X(_11699_));
 sky130_fd_sc_hd__o32a_2 _15238_ (.A1(instr_jalr),
    .A2(_10723_),
    .A3(_11697_),
    .B1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B2(_11699_),
    .X(_03207_));
 sky130_fd_sc_hd__buf_1 _15239_ (.A(is_slli_srli_srai),
    .X(_11700_));
 sky130_fd_sc_hd__buf_1 _15240_ (.A(_10760_),
    .X(_11701_));
 sky130_fd_sc_hd__o31a_2 _15241_ (.A1(_10740_),
    .A2(_00334_),
    .A3(_10744_),
    .B1(_10732_),
    .X(_11702_));
 sky130_fd_sc_hd__or4_2 _15242_ (.A(_10738_),
    .B(_10726_),
    .C(_10768_),
    .D(_10722_),
    .X(_11703_));
 sky130_fd_sc_hd__o2bb2ai_2 _15243_ (.A1_N(_11700_),
    .A2_N(_11701_),
    .B1(_11702_),
    .B2(_11703_),
    .Y(_03206_));
 sky130_fd_sc_hd__o32a_2 _15244_ (.A1(_00329_),
    .A2(_10714_),
    .A3(_11647_),
    .B1(_10663_),
    .B2(_10493_),
    .X(_11704_));
 sky130_vsdinv _15245_ (.A(_11704_),
    .Y(_03205_));
 sky130_fd_sc_hd__buf_1 _15246_ (.A(\decoded_imm_uj[20] ),
    .X(_11705_));
 sky130_fd_sc_hd__buf_1 _15247_ (.A(_11705_),
    .X(_11706_));
 sky130_fd_sc_hd__buf_1 _15248_ (.A(_11706_),
    .X(_11707_));
 sky130_fd_sc_hd__buf_1 _15249_ (.A(_10718_),
    .X(_11708_));
 sky130_fd_sc_hd__a22o_2 _15250_ (.A1(_11707_),
    .A2(_11708_),
    .B1(\mem_rdata_latched[31] ),
    .B2(_12947_),
    .X(_03204_));
 sky130_fd_sc_hd__a22o_2 _15251_ (.A1(\decoded_imm_uj[19] ),
    .A2(_11708_),
    .B1(\mem_rdata_latched[19] ),
    .B2(_12947_),
    .X(_03203_));
 sky130_fd_sc_hd__buf_1 _15252_ (.A(_10492_),
    .X(_11709_));
 sky130_fd_sc_hd__buf_1 _15253_ (.A(_10718_),
    .X(_11710_));
 sky130_fd_sc_hd__a22o_2 _15254_ (.A1(\mem_rdata_latched[18] ),
    .A2(_11709_),
    .B1(\decoded_imm_uj[18] ),
    .B2(_11710_),
    .X(_03202_));
 sky130_fd_sc_hd__a22o_2 _15255_ (.A1(\mem_rdata_latched[17] ),
    .A2(_10717_),
    .B1(\decoded_imm_uj[17] ),
    .B2(_11710_),
    .X(_03201_));
 sky130_fd_sc_hd__a22o_2 _15256_ (.A1(\mem_rdata_latched[16] ),
    .A2(_10717_),
    .B1(\decoded_imm_uj[16] ),
    .B2(_11710_),
    .X(_03200_));
 sky130_fd_sc_hd__a22o_2 _15257_ (.A1(\mem_rdata_latched[15] ),
    .A2(_10717_),
    .B1(\decoded_imm_uj[15] ),
    .B2(_11710_),
    .X(_03199_));
 sky130_fd_sc_hd__a22o_2 _15258_ (.A1(\decoded_imm_uj[14] ),
    .A2(_11708_),
    .B1(\mem_rdata_latched[14] ),
    .B2(_12947_),
    .X(_03198_));
 sky130_fd_sc_hd__buf_1 _15259_ (.A(_10493_),
    .X(_11711_));
 sky130_fd_sc_hd__a22o_2 _15260_ (.A1(\decoded_imm_uj[13] ),
    .A2(_11708_),
    .B1(\mem_rdata_latched[13] ),
    .B2(_11711_),
    .X(_03197_));
 sky130_fd_sc_hd__a22o_2 _15261_ (.A1(\decoded_imm_uj[12] ),
    .A2(_11708_),
    .B1(\mem_rdata_latched[12] ),
    .B2(_11711_),
    .X(_03196_));
 sky130_fd_sc_hd__a22o_2 _15262_ (.A1(\decoded_imm_uj[11] ),
    .A2(_11708_),
    .B1(\mem_rdata_latched[20] ),
    .B2(_11711_),
    .X(_03195_));
 sky130_fd_sc_hd__buf_1 _15263_ (.A(_10718_),
    .X(_11712_));
 sky130_fd_sc_hd__a22o_2 _15264_ (.A1(\decoded_imm_uj[10] ),
    .A2(_11712_),
    .B1(\mem_rdata_latched[30] ),
    .B2(_11711_),
    .X(_03194_));
 sky130_fd_sc_hd__a22o_2 _15265_ (.A1(\decoded_imm_uj[9] ),
    .A2(_11712_),
    .B1(\mem_rdata_latched[29] ),
    .B2(_11711_),
    .X(_03193_));
 sky130_fd_sc_hd__a22o_2 _15266_ (.A1(\decoded_imm_uj[8] ),
    .A2(_11712_),
    .B1(\mem_rdata_latched[28] ),
    .B2(_11711_),
    .X(_03192_));
 sky130_fd_sc_hd__a22o_2 _15267_ (.A1(\mem_rdata_latched[27] ),
    .A2(_10717_),
    .B1(\decoded_imm_uj[7] ),
    .B2(_11710_),
    .X(_03191_));
 sky130_fd_sc_hd__buf_1 _15268_ (.A(_10492_),
    .X(_11713_));
 sky130_fd_sc_hd__a22o_2 _15269_ (.A1(\decoded_imm_uj[6] ),
    .A2(_11712_),
    .B1(\mem_rdata_latched[26] ),
    .B2(_11713_),
    .X(_03190_));
 sky130_fd_sc_hd__a22o_2 _15270_ (.A1(\decoded_imm_uj[5] ),
    .A2(_11712_),
    .B1(\mem_rdata_latched[25] ),
    .B2(_11713_),
    .X(_03189_));
 sky130_fd_sc_hd__a22o_2 _15271_ (.A1(\decoded_imm_uj[4] ),
    .A2(_11712_),
    .B1(\mem_rdata_latched[24] ),
    .B2(_11713_),
    .X(_03188_));
 sky130_fd_sc_hd__buf_1 _15272_ (.A(_10718_),
    .X(_11714_));
 sky130_fd_sc_hd__a22o_2 _15273_ (.A1(\decoded_imm_uj[3] ),
    .A2(_11714_),
    .B1(\mem_rdata_latched[23] ),
    .B2(_11713_),
    .X(_03187_));
 sky130_fd_sc_hd__a22o_2 _15274_ (.A1(\decoded_imm_uj[2] ),
    .A2(_11714_),
    .B1(\mem_rdata_latched[22] ),
    .B2(_11713_),
    .X(_03186_));
 sky130_fd_sc_hd__a22o_2 _15275_ (.A1(\decoded_imm_uj[1] ),
    .A2(_11714_),
    .B1(\mem_rdata_latched[21] ),
    .B2(_11713_),
    .X(_03185_));
 sky130_fd_sc_hd__inv_2 _15276_ (.A(\decoded_imm[0] ),
    .Y(_11715_));
 sky130_fd_sc_hd__buf_1 _15277_ (.A(_11698_),
    .X(_11716_));
 sky130_vsdinv _15278_ (.A(\mem_rdata_q[7] ),
    .Y(_11717_));
 sky130_vsdinv _15279_ (.A(\mem_rdata_q[20] ),
    .Y(_11718_));
 sky130_fd_sc_hd__or3_2 _15280_ (.A(is_alu_reg_imm),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(instr_jalr),
    .X(_11719_));
 sky130_vsdinv _15281_ (.A(_11719_),
    .Y(_11720_));
 sky130_fd_sc_hd__o22a_2 _15282_ (.A1(_10666_),
    .A2(_11717_),
    .B1(_11718_),
    .B2(_11720_),
    .X(_11721_));
 sky130_fd_sc_hd__o22ai_2 _15283_ (.A1(_11715_),
    .A2(_11716_),
    .B1(_11701_),
    .B2(_11721_),
    .Y(_03184_));
 sky130_fd_sc_hd__a22o_2 _15284_ (.A1(\decoded_rd[4] ),
    .A2(_11714_),
    .B1(\mem_rdata_latched[11] ),
    .B2(_11709_),
    .X(_03183_));
 sky130_fd_sc_hd__a22o_2 _15285_ (.A1(\decoded_rd[3] ),
    .A2(_11714_),
    .B1(\mem_rdata_latched[10] ),
    .B2(_11709_),
    .X(_03182_));
 sky130_fd_sc_hd__a22o_2 _15286_ (.A1(\decoded_rd[2] ),
    .A2(_11714_),
    .B1(\mem_rdata_latched[9] ),
    .B2(_11709_),
    .X(_03181_));
 sky130_fd_sc_hd__a22o_2 _15287_ (.A1(\decoded_rd[1] ),
    .A2(_10494_),
    .B1(\mem_rdata_latched[8] ),
    .B2(_11709_),
    .X(_03180_));
 sky130_fd_sc_hd__a22o_2 _15288_ (.A1(\decoded_rd[0] ),
    .A2(_10494_),
    .B1(\mem_rdata_latched[7] ),
    .B2(_11709_),
    .X(_03179_));
 sky130_fd_sc_hd__buf_1 _15289_ (.A(\mem_rdata_q[27] ),
    .X(_11722_));
 sky130_vsdinv _15290_ (.A(_11722_),
    .Y(_11723_));
 sky130_fd_sc_hd__or2_2 _15291_ (.A(_11723_),
    .B(_10741_),
    .X(_11724_));
 sky130_vsdinv _15292_ (.A(\mem_rdata_q[1] ),
    .Y(_11725_));
 sky130_vsdinv _15293_ (.A(\mem_rdata_q[0] ),
    .Y(_11726_));
 sky130_fd_sc_hd__or4_2 _15294_ (.A(_11725_),
    .B(_11726_),
    .C(\mem_rdata_q[6] ),
    .D(\mem_rdata_q[5] ),
    .X(_11727_));
 sky130_fd_sc_hd__or4b_2 _15295_ (.A(\mem_rdata_q[4] ),
    .B(_11727_),
    .C(\mem_rdata_q[2] ),
    .D_N(\mem_rdata_q[3] ),
    .X(_11728_));
 sky130_fd_sc_hd__buf_1 _15296_ (.A(\mem_rdata_q[28] ),
    .X(_11729_));
 sky130_fd_sc_hd__buf_1 _15297_ (.A(\mem_rdata_q[26] ),
    .X(_11730_));
 sky130_vsdinv _15298_ (.A(\mem_rdata_q[25] ),
    .Y(_11731_));
 sky130_fd_sc_hd__or4_2 _15299_ (.A(_10742_),
    .B(\mem_rdata_q[30] ),
    .C(\mem_rdata_q[29] ),
    .D(_11731_),
    .X(_11732_));
 sky130_fd_sc_hd__or3_2 _15300_ (.A(_11729_),
    .B(_11730_),
    .C(_11732_),
    .X(_11733_));
 sky130_vsdinv _15301_ (.A(instr_timer),
    .Y(_11734_));
 sky130_fd_sc_hd__buf_1 _15302_ (.A(_11734_),
    .X(_11735_));
 sky130_fd_sc_hd__buf_1 _15303_ (.A(_10748_),
    .X(_11736_));
 sky130_fd_sc_hd__o32a_2 _15304_ (.A1(_11724_),
    .A2(_11728_),
    .A3(_11733_),
    .B1(_11735_),
    .B2(_11736_),
    .X(_11737_));
 sky130_vsdinv _15305_ (.A(_11737_),
    .Y(_03178_));
 sky130_fd_sc_hd__nor2_2 _15306_ (.A(_10500_),
    .B(_10503_),
    .Y(_11738_));
 sky130_fd_sc_hd__a32o_2 _15307_ (.A1(\mem_rdata_latched[27] ),
    .A2(_10506_),
    .A3(_11738_),
    .B1(instr_waitirq),
    .B2(_10719_),
    .X(_03177_));
 sky130_vsdinv _15308_ (.A(_11730_),
    .Y(_11739_));
 sky130_fd_sc_hd__or4_2 _15309_ (.A(_11739_),
    .B(_10721_),
    .C(_11729_),
    .D(_11722_),
    .X(_11740_));
 sky130_fd_sc_hd__buf_1 _15310_ (.A(_10678_),
    .X(_11741_));
 sky130_fd_sc_hd__o32a_2 _15311_ (.A1(_11732_),
    .A2(_11740_),
    .A3(_11728_),
    .B1(_11741_),
    .B2(_11736_),
    .X(_11742_));
 sky130_vsdinv _15312_ (.A(_11742_),
    .Y(_03176_));
 sky130_fd_sc_hd__a2bb2o_2 _15313_ (.A1_N(_00337_),
    .A2_N(_10505_),
    .B1(instr_retirq),
    .B2(_00337_),
    .X(_03175_));
 sky130_fd_sc_hd__buf_1 _15314_ (.A(_10749_),
    .X(_11743_));
 sky130_fd_sc_hd__or4_2 _15315_ (.A(_11722_),
    .B(_10722_),
    .C(_11728_),
    .D(_11733_),
    .X(_11744_));
 sky130_fd_sc_hd__o21ai_2 _15316_ (.A1(_11425_),
    .A2(_11743_),
    .B1(_11744_),
    .Y(_03174_));
 sky130_fd_sc_hd__buf_1 _15317_ (.A(_10741_),
    .X(_11745_));
 sky130_fd_sc_hd__buf_1 _15318_ (.A(_11745_),
    .X(_11746_));
 sky130_vsdinv _15319_ (.A(_10733_),
    .Y(_11747_));
 sky130_vsdinv _15320_ (.A(_11728_),
    .Y(_11748_));
 sky130_fd_sc_hd__a22o_2 _15321_ (.A1(instr_getq),
    .A2(_11746_),
    .B1(_11747_),
    .B2(_11748_),
    .X(_03173_));
 sky130_fd_sc_hd__or2_2 _15322_ (.A(\mem_rdata_q[23] ),
    .B(\mem_rdata_q[22] ),
    .X(_11749_));
 sky130_fd_sc_hd__or4_2 _15323_ (.A(\mem_rdata_q[11] ),
    .B(\mem_rdata_q[10] ),
    .C(\mem_rdata_q[8] ),
    .D(\mem_rdata_q[7] ),
    .X(_11750_));
 sky130_fd_sc_hd__or4_2 _15324_ (.A(\mem_rdata_q[24] ),
    .B(\mem_rdata_q[21] ),
    .C(_11749_),
    .D(_11750_),
    .X(_11751_));
 sky130_fd_sc_hd__or4_2 _15325_ (.A(\mem_rdata_q[9] ),
    .B(_10722_),
    .C(_10763_),
    .D(_11751_),
    .X(_11752_));
 sky130_fd_sc_hd__or2_2 _15326_ (.A(\mem_rdata_q[19] ),
    .B(\mem_rdata_q[18] ),
    .X(_11753_));
 sky130_fd_sc_hd__or4_2 _15327_ (.A(\mem_rdata_q[17] ),
    .B(\mem_rdata_q[16] ),
    .C(\mem_rdata_q[15] ),
    .D(_11753_),
    .X(_11754_));
 sky130_fd_sc_hd__or4bb_2 _15328_ (.A(_11725_),
    .B(_11726_),
    .C_N(\mem_rdata_q[6] ),
    .D_N(\mem_rdata_q[5] ),
    .X(_11755_));
 sky130_fd_sc_hd__or4b_2 _15329_ (.A(_11755_),
    .B(\mem_rdata_q[3] ),
    .C(\mem_rdata_q[2] ),
    .D_N(\mem_rdata_q[4] ),
    .X(_11756_));
 sky130_fd_sc_hd__or3_2 _15330_ (.A(_10732_),
    .B(_11754_),
    .C(_11756_),
    .X(_11757_));
 sky130_fd_sc_hd__o2bb2ai_2 _15331_ (.A1_N(instr_ecall_ebreak),
    .A2_N(_11701_),
    .B1(_11752_),
    .B2(_11757_),
    .Y(_03172_));
 sky130_vsdinv _15332_ (.A(\mem_rdata_q[21] ),
    .Y(_11758_));
 sky130_fd_sc_hd__or2_2 _15333_ (.A(_11758_),
    .B(_11749_),
    .X(_11759_));
 sky130_fd_sc_hd__or4_2 _15334_ (.A(\mem_rdata_q[20] ),
    .B(_10721_),
    .C(_11759_),
    .D(_11756_),
    .X(_11760_));
 sky130_vsdinv _15335_ (.A(_10742_),
    .Y(_11761_));
 sky130_fd_sc_hd__or4_2 _15336_ (.A(_11761_),
    .B(_10743_),
    .C(_10740_),
    .D(_11729_),
    .X(_11762_));
 sky130_fd_sc_hd__or2_2 _15337_ (.A(\mem_rdata_q[25] ),
    .B(\mem_rdata_q[24] ),
    .X(_11763_));
 sky130_fd_sc_hd__or4_2 _15338_ (.A(_11762_),
    .B(_11763_),
    .C(_11723_),
    .D(_11730_),
    .X(_11764_));
 sky130_fd_sc_hd__or2_2 _15339_ (.A(_10758_),
    .B(_11754_),
    .X(_11765_));
 sky130_fd_sc_hd__buf_1 _15340_ (.A(_10616_),
    .X(_11766_));
 sky130_fd_sc_hd__o32a_2 _15341_ (.A1(_11760_),
    .A2(_11764_),
    .A3(_11765_),
    .B1(_11766_),
    .B2(_11736_),
    .X(_11767_));
 sky130_vsdinv _15342_ (.A(_11767_),
    .Y(_03171_));
 sky130_fd_sc_hd__buf_1 _15343_ (.A(_10617_),
    .X(_11768_));
 sky130_fd_sc_hd__or3_2 _15344_ (.A(\mem_rdata_q[29] ),
    .B(\mem_rdata_q[28] ),
    .C(\mem_rdata_q[25] ),
    .X(_11769_));
 sky130_fd_sc_hd__or4_2 _15345_ (.A(_11761_),
    .B(_10743_),
    .C(_11769_),
    .D(_11722_),
    .X(_11770_));
 sky130_fd_sc_hd__or4_2 _15346_ (.A(_11730_),
    .B(\mem_rdata_q[24] ),
    .C(_11765_),
    .D(_11770_),
    .X(_11771_));
 sky130_fd_sc_hd__o22ai_2 _15347_ (.A1(_11768_),
    .A2(_11716_),
    .B1(_11760_),
    .B2(_11771_),
    .Y(_03170_));
 sky130_fd_sc_hd__or4_2 _15348_ (.A(\mem_rdata_q[21] ),
    .B(_10721_),
    .C(_11749_),
    .D(_11756_),
    .X(_11772_));
 sky130_fd_sc_hd__buf_1 _15349_ (.A(_10618_),
    .X(_11773_));
 sky130_fd_sc_hd__o32a_2 _15350_ (.A1(_11764_),
    .A2(_11772_),
    .A3(_11765_),
    .B1(_11773_),
    .B2(_11736_),
    .X(_11774_));
 sky130_vsdinv _15351_ (.A(_11774_),
    .Y(_03169_));
 sky130_fd_sc_hd__o22ai_2 _15352_ (.A1(_10615_),
    .A2(_11716_),
    .B1(_11771_),
    .B2(_11772_),
    .Y(_03168_));
 sky130_vsdinv _15353_ (.A(_10739_),
    .Y(_11775_));
 sky130_vsdinv _15354_ (.A(_10745_),
    .Y(_11776_));
 sky130_fd_sc_hd__buf_1 _15355_ (.A(_10760_),
    .X(_11777_));
 sky130_fd_sc_hd__a32o_2 _15356_ (.A1(is_alu_reg_imm),
    .A2(_11775_),
    .A3(_11776_),
    .B1(instr_srai),
    .B2(_11777_),
    .X(_03167_));
 sky130_fd_sc_hd__a32o_2 _15357_ (.A1(is_alu_reg_imm),
    .A2(_11775_),
    .A3(_11747_),
    .B1(instr_srli),
    .B2(_11777_),
    .X(_03166_));
 sky130_vsdinv _15358_ (.A(_10761_),
    .Y(_11778_));
 sky130_fd_sc_hd__a32o_2 _15359_ (.A1(is_alu_reg_imm),
    .A2(_11778_),
    .A3(_11747_),
    .B1(instr_slli),
    .B2(_11777_),
    .X(_03165_));
 sky130_vsdinv _15360_ (.A(instr_sw),
    .Y(_11779_));
 sky130_fd_sc_hd__o32a_2 _15361_ (.A1(_10666_),
    .A2(_10722_),
    .A3(_10758_),
    .B1(_11779_),
    .B2(_11736_),
    .X(_11780_));
 sky130_vsdinv _15362_ (.A(_11780_),
    .Y(_03164_));
 sky130_fd_sc_hd__buf_1 _15363_ (.A(_10747_),
    .X(_11781_));
 sky130_fd_sc_hd__buf_1 _15364_ (.A(_11781_),
    .X(_11782_));
 sky130_fd_sc_hd__a32o_2 _15365_ (.A1(_10665_),
    .A2(_11782_),
    .A3(_11778_),
    .B1(instr_sh),
    .B2(_11777_),
    .X(_03163_));
 sky130_vsdinv _15366_ (.A(_10763_),
    .Y(_11783_));
 sky130_fd_sc_hd__a32o_2 _15367_ (.A1(_10665_),
    .A2(_11782_),
    .A3(_11783_),
    .B1(instr_sb),
    .B2(_11777_),
    .X(_03162_));
 sky130_fd_sc_hd__a32o_2 _15368_ (.A1(is_lb_lh_lw_lbu_lhu),
    .A2(_11782_),
    .A3(_11775_),
    .B1(instr_lhu),
    .B2(_11777_),
    .X(_03161_));
 sky130_vsdinv _15369_ (.A(_10753_),
    .Y(_11784_));
 sky130_fd_sc_hd__buf_1 _15370_ (.A(_11745_),
    .X(_11785_));
 sky130_fd_sc_hd__a32o_2 _15371_ (.A1(is_lb_lh_lw_lbu_lhu),
    .A2(_11782_),
    .A3(_11784_),
    .B1(instr_lbu),
    .B2(_11785_),
    .X(_03160_));
 sky130_vsdinv _15372_ (.A(instr_lw),
    .Y(_11786_));
 sky130_fd_sc_hd__o32a_2 _15373_ (.A1(_10663_),
    .A2(_10722_),
    .A3(_10758_),
    .B1(_11786_),
    .B2(_11736_),
    .X(_11787_));
 sky130_vsdinv _15374_ (.A(_11787_),
    .Y(_03159_));
 sky130_fd_sc_hd__buf_1 _15375_ (.A(_11781_),
    .X(_11788_));
 sky130_fd_sc_hd__a32o_2 _15376_ (.A1(is_lb_lh_lw_lbu_lhu),
    .A2(_11788_),
    .A3(_11778_),
    .B1(instr_lh),
    .B2(_11785_),
    .X(_03158_));
 sky130_fd_sc_hd__a32o_2 _15377_ (.A1(is_lb_lh_lw_lbu_lhu),
    .A2(_11788_),
    .A3(_11783_),
    .B1(instr_lb),
    .B2(_11785_),
    .X(_03157_));
 sky130_fd_sc_hd__or3b_2 _15378_ (.A(_10497_),
    .B(_10498_),
    .C_N(_00326_),
    .X(_11789_));
 sky130_fd_sc_hd__or2_2 _15379_ (.A(_00327_),
    .B(_11789_),
    .X(_11790_));
 sky130_fd_sc_hd__or4_2 _15380_ (.A(\mem_rdata_latched[14] ),
    .B(\mem_rdata_latched[13] ),
    .C(\mem_rdata_latched[12] ),
    .D(_10715_),
    .X(_11791_));
 sky130_vsdinv _15381_ (.A(instr_jalr),
    .Y(_02063_));
 sky130_fd_sc_hd__o32a_2 _15382_ (.A1(_11790_),
    .A2(_11791_),
    .A3(_10718_),
    .B1(_02063_),
    .B2(_10493_),
    .X(_11792_));
 sky130_vsdinv _15383_ (.A(_11792_),
    .Y(_03156_));
 sky130_vsdinv _15384_ (.A(instr_jal),
    .Y(_11793_));
 sky130_fd_sc_hd__buf_1 _15385_ (.A(_11793_),
    .X(_11794_));
 sky130_fd_sc_hd__buf_1 _15386_ (.A(_11794_),
    .X(_00323_));
 sky130_fd_sc_hd__or3_2 _15387_ (.A(_10495_),
    .B(_10715_),
    .C(_11789_),
    .X(_11795_));
 sky130_fd_sc_hd__o22ai_2 _15388_ (.A1(_00323_),
    .A2(_12947_),
    .B1(_00337_),
    .B2(_11795_),
    .Y(_03155_));
 sky130_fd_sc_hd__nor3_2 _15389_ (.A(_00330_),
    .B(_10494_),
    .C(_11790_),
    .Y(_11796_));
 sky130_fd_sc_hd__a32o_2 _15390_ (.A1(_10713_),
    .A2(_10714_),
    .A3(_11796_),
    .B1(instr_auipc),
    .B2(_10719_),
    .X(_03154_));
 sky130_fd_sc_hd__buf_1 _15391_ (.A(instr_lui),
    .X(_11797_));
 sky130_fd_sc_hd__a32o_2 _15392_ (.A1(_00329_),
    .A2(_10714_),
    .A3(_11796_),
    .B1(_11797_),
    .B2(_11710_),
    .X(_03153_));
 sky130_fd_sc_hd__buf_1 _15393_ (.A(_11698_),
    .X(_11798_));
 sky130_fd_sc_hd__a22o_2 _15394_ (.A1(pcpi_insn[31]),
    .A2(_11746_),
    .B1(_10742_),
    .B2(_11798_),
    .X(_03152_));
 sky130_fd_sc_hd__buf_1 _15395_ (.A(_11781_),
    .X(_11799_));
 sky130_fd_sc_hd__a22o_2 _15396_ (.A1(pcpi_insn[30]),
    .A2(_11746_),
    .B1(\mem_rdata_q[30] ),
    .B2(_11799_),
    .X(_03151_));
 sky130_fd_sc_hd__o22a_2 _15397_ (.A1(_10740_),
    .A2(_11785_),
    .B1(pcpi_insn[29]),
    .B2(_11743_),
    .X(_03150_));
 sky130_fd_sc_hd__buf_1 _15398_ (.A(_11745_),
    .X(_11800_));
 sky130_fd_sc_hd__a22o_2 _15399_ (.A1(pcpi_insn[28]),
    .A2(_11800_),
    .B1(_11729_),
    .B2(_11799_),
    .X(_03149_));
 sky130_fd_sc_hd__o22a_2 _15400_ (.A1(_11722_),
    .A2(_11785_),
    .B1(pcpi_insn[27]),
    .B2(_11743_),
    .X(_03148_));
 sky130_fd_sc_hd__a22o_2 _15401_ (.A1(_11730_),
    .A2(_11782_),
    .B1(pcpi_insn[26]),
    .B2(_11785_),
    .X(_03147_));
 sky130_fd_sc_hd__a22o_2 _15402_ (.A1(pcpi_insn[25]),
    .A2(_11800_),
    .B1(\mem_rdata_q[25] ),
    .B2(_11799_),
    .X(_03146_));
 sky130_fd_sc_hd__a22o_2 _15403_ (.A1(pcpi_insn[24]),
    .A2(_11800_),
    .B1(\mem_rdata_q[24] ),
    .B2(_11799_),
    .X(_03145_));
 sky130_fd_sc_hd__a22o_2 _15404_ (.A1(pcpi_insn[23]),
    .A2(_11800_),
    .B1(\mem_rdata_q[23] ),
    .B2(_11799_),
    .X(_03144_));
 sky130_fd_sc_hd__a22o_2 _15405_ (.A1(pcpi_insn[22]),
    .A2(_11800_),
    .B1(\mem_rdata_q[22] ),
    .B2(_11799_),
    .X(_03143_));
 sky130_fd_sc_hd__o22a_2 _15406_ (.A1(\mem_rdata_q[21] ),
    .A2(_11746_),
    .B1(pcpi_insn[21]),
    .B2(_11743_),
    .X(_03142_));
 sky130_fd_sc_hd__o22a_2 _15407_ (.A1(\mem_rdata_q[20] ),
    .A2(_11746_),
    .B1(pcpi_insn[20]),
    .B2(_11743_),
    .X(_03141_));
 sky130_fd_sc_hd__buf_1 _15408_ (.A(_11781_),
    .X(_11801_));
 sky130_fd_sc_hd__a22o_2 _15409_ (.A1(pcpi_insn[19]),
    .A2(_11800_),
    .B1(\mem_rdata_q[19] ),
    .B2(_11801_),
    .X(_03140_));
 sky130_fd_sc_hd__buf_1 _15410_ (.A(_11745_),
    .X(_11802_));
 sky130_fd_sc_hd__a22o_2 _15411_ (.A1(pcpi_insn[18]),
    .A2(_11802_),
    .B1(\mem_rdata_q[18] ),
    .B2(_11801_),
    .X(_03139_));
 sky130_fd_sc_hd__a22o_2 _15412_ (.A1(pcpi_insn[17]),
    .A2(_11802_),
    .B1(\mem_rdata_q[17] ),
    .B2(_11801_),
    .X(_03138_));
 sky130_fd_sc_hd__a22o_2 _15413_ (.A1(pcpi_insn[16]),
    .A2(_11802_),
    .B1(\mem_rdata_q[16] ),
    .B2(_11801_),
    .X(_03137_));
 sky130_fd_sc_hd__a22o_2 _15414_ (.A1(pcpi_insn[15]),
    .A2(_11802_),
    .B1(\mem_rdata_q[15] ),
    .B2(_11801_),
    .X(_03136_));
 sky130_fd_sc_hd__a22o_2 _15415_ (.A1(pcpi_insn[14]),
    .A2(_11802_),
    .B1(_10727_),
    .B2(_11801_),
    .X(_03135_));
 sky130_fd_sc_hd__buf_1 _15416_ (.A(_11781_),
    .X(_11803_));
 sky130_fd_sc_hd__a22o_2 _15417_ (.A1(pcpi_insn[13]),
    .A2(_11802_),
    .B1(_10738_),
    .B2(_11803_),
    .X(_03134_));
 sky130_fd_sc_hd__buf_1 _15418_ (.A(_11745_),
    .X(_11804_));
 sky130_fd_sc_hd__a22o_2 _15419_ (.A1(pcpi_insn[12]),
    .A2(_11804_),
    .B1(_10725_),
    .B2(_11803_),
    .X(_03133_));
 sky130_fd_sc_hd__a22o_2 _15420_ (.A1(pcpi_insn[11]),
    .A2(_11804_),
    .B1(\mem_rdata_q[11] ),
    .B2(_11803_),
    .X(_03132_));
 sky130_fd_sc_hd__a22o_2 _15421_ (.A1(pcpi_insn[10]),
    .A2(_11804_),
    .B1(\mem_rdata_q[10] ),
    .B2(_11803_),
    .X(_03131_));
 sky130_fd_sc_hd__o22a_2 _15422_ (.A1(\mem_rdata_q[9] ),
    .A2(_11746_),
    .B1(pcpi_insn[9]),
    .B2(_11743_),
    .X(_03130_));
 sky130_fd_sc_hd__a22o_2 _15423_ (.A1(pcpi_insn[8]),
    .A2(_11804_),
    .B1(\mem_rdata_q[8] ),
    .B2(_11803_),
    .X(_03129_));
 sky130_fd_sc_hd__a22o_2 _15424_ (.A1(pcpi_insn[7]),
    .A2(_11804_),
    .B1(\mem_rdata_q[7] ),
    .B2(_11803_),
    .X(_03128_));
 sky130_fd_sc_hd__buf_1 _15425_ (.A(_11781_),
    .X(_11805_));
 sky130_fd_sc_hd__a22o_2 _15426_ (.A1(pcpi_insn[6]),
    .A2(_11804_),
    .B1(\mem_rdata_q[6] ),
    .B2(_11805_),
    .X(_03127_));
 sky130_fd_sc_hd__buf_1 _15427_ (.A(_11745_),
    .X(_11806_));
 sky130_fd_sc_hd__a22o_2 _15428_ (.A1(pcpi_insn[5]),
    .A2(_11806_),
    .B1(\mem_rdata_q[5] ),
    .B2(_11805_),
    .X(_03126_));
 sky130_fd_sc_hd__a22o_2 _15429_ (.A1(pcpi_insn[4]),
    .A2(_11806_),
    .B1(\mem_rdata_q[4] ),
    .B2(_11805_),
    .X(_03125_));
 sky130_fd_sc_hd__a22o_2 _15430_ (.A1(pcpi_insn[3]),
    .A2(_11806_),
    .B1(\mem_rdata_q[3] ),
    .B2(_11805_),
    .X(_03124_));
 sky130_fd_sc_hd__a22o_2 _15431_ (.A1(pcpi_insn[2]),
    .A2(_11806_),
    .B1(\mem_rdata_q[2] ),
    .B2(_11805_),
    .X(_03123_));
 sky130_fd_sc_hd__a22o_2 _15432_ (.A1(pcpi_insn[1]),
    .A2(_11806_),
    .B1(\mem_rdata_q[1] ),
    .B2(_11805_),
    .X(_03122_));
 sky130_fd_sc_hd__a22o_2 _15433_ (.A1(pcpi_insn[0]),
    .A2(_11806_),
    .B1(\mem_rdata_q[0] ),
    .B2(_11782_),
    .X(_03121_));
 sky130_vsdinv _15434_ (.A(\cpu_state[5] ),
    .Y(_11807_));
 sky130_fd_sc_hd__and3_2 _15435_ (.A(_10468_),
    .B(_10458_),
    .C(_11807_),
    .X(_11808_));
 sky130_fd_sc_hd__or4_2 _15436_ (.A(_10476_),
    .B(_00318_),
    .C(_00320_),
    .D(_11808_),
    .X(_11809_));
 sky130_fd_sc_hd__buf_1 _15437_ (.A(_11809_),
    .X(_11810_));
 sky130_fd_sc_hd__buf_1 _15438_ (.A(_11810_),
    .X(_11811_));
 sky130_fd_sc_hd__buf_1 _15439_ (.A(pcpi_rs1[31]),
    .X(_11812_));
 sky130_vsdinv _15440_ (.A(_11809_),
    .Y(_11813_));
 sky130_fd_sc_hd__buf_1 _15441_ (.A(_11813_),
    .X(_11814_));
 sky130_fd_sc_hd__buf_1 _15442_ (.A(_11814_),
    .X(_11815_));
 sky130_fd_sc_hd__o22a_2 _15443_ (.A1(_02499_),
    .A2(_11811_),
    .B1(_11812_),
    .B2(_11815_),
    .X(_03120_));
 sky130_fd_sc_hd__buf_1 _15444_ (.A(pcpi_rs1[30]),
    .X(_11816_));
 sky130_fd_sc_hd__o22a_2 _15445_ (.A1(_02498_),
    .A2(_11811_),
    .B1(_11816_),
    .B2(_11815_),
    .X(_03119_));
 sky130_fd_sc_hd__buf_1 _15446_ (.A(pcpi_rs1[29]),
    .X(_11817_));
 sky130_fd_sc_hd__o22a_2 _15447_ (.A1(_02496_),
    .A2(_11811_),
    .B1(_11817_),
    .B2(_11815_),
    .X(_03118_));
 sky130_fd_sc_hd__buf_1 _15448_ (.A(pcpi_rs1[28]),
    .X(_11818_));
 sky130_fd_sc_hd__o22a_2 _15449_ (.A1(_02495_),
    .A2(_11811_),
    .B1(_11818_),
    .B2(_11815_),
    .X(_03117_));
 sky130_fd_sc_hd__buf_1 _15450_ (.A(pcpi_rs1[27]),
    .X(_11819_));
 sky130_fd_sc_hd__buf_1 _15451_ (.A(_11819_),
    .X(_11820_));
 sky130_fd_sc_hd__o22a_2 _15452_ (.A1(_02494_),
    .A2(_11811_),
    .B1(_11820_),
    .B2(_11815_),
    .X(_03116_));
 sky130_fd_sc_hd__buf_1 _15453_ (.A(pcpi_rs1[26]),
    .X(_11821_));
 sky130_fd_sc_hd__buf_1 _15454_ (.A(_11821_),
    .X(_11822_));
 sky130_fd_sc_hd__o22a_2 _15455_ (.A1(_02493_),
    .A2(_11811_),
    .B1(_11822_),
    .B2(_11815_),
    .X(_03115_));
 sky130_fd_sc_hd__buf_1 _15456_ (.A(_11810_),
    .X(_11823_));
 sky130_fd_sc_hd__buf_1 _15457_ (.A(pcpi_rs1[25]),
    .X(_11824_));
 sky130_fd_sc_hd__buf_1 _15458_ (.A(_11824_),
    .X(_11825_));
 sky130_fd_sc_hd__buf_1 _15459_ (.A(_11814_),
    .X(_11826_));
 sky130_fd_sc_hd__o22a_2 _15460_ (.A1(_02492_),
    .A2(_11823_),
    .B1(_11825_),
    .B2(_11826_),
    .X(_03114_));
 sky130_fd_sc_hd__buf_1 _15461_ (.A(pcpi_rs1[24]),
    .X(_11827_));
 sky130_fd_sc_hd__buf_1 _15462_ (.A(_11827_),
    .X(_11828_));
 sky130_fd_sc_hd__o22a_2 _15463_ (.A1(_02491_),
    .A2(_11823_),
    .B1(_11828_),
    .B2(_11826_),
    .X(_03113_));
 sky130_fd_sc_hd__buf_1 _15464_ (.A(pcpi_rs1[23]),
    .X(_11829_));
 sky130_fd_sc_hd__o22a_2 _15465_ (.A1(_02490_),
    .A2(_11823_),
    .B1(_11829_),
    .B2(_11826_),
    .X(_03112_));
 sky130_fd_sc_hd__buf_1 _15466_ (.A(pcpi_rs1[22]),
    .X(_11830_));
 sky130_fd_sc_hd__o22a_2 _15467_ (.A1(_02489_),
    .A2(_11823_),
    .B1(_11830_),
    .B2(_11826_),
    .X(_03111_));
 sky130_fd_sc_hd__buf_1 _15468_ (.A(pcpi_rs1[21]),
    .X(_11831_));
 sky130_fd_sc_hd__o22a_2 _15469_ (.A1(_02488_),
    .A2(_11823_),
    .B1(_11831_),
    .B2(_11826_),
    .X(_03110_));
 sky130_fd_sc_hd__buf_1 _15470_ (.A(pcpi_rs1[20]),
    .X(_11832_));
 sky130_fd_sc_hd__o22a_2 _15471_ (.A1(_02487_),
    .A2(_11823_),
    .B1(_11832_),
    .B2(_11826_),
    .X(_03109_));
 sky130_fd_sc_hd__buf_1 _15472_ (.A(_11810_),
    .X(_11833_));
 sky130_fd_sc_hd__buf_1 _15473_ (.A(pcpi_rs1[19]),
    .X(_11834_));
 sky130_fd_sc_hd__buf_1 _15474_ (.A(_11814_),
    .X(_11835_));
 sky130_fd_sc_hd__o22a_2 _15475_ (.A1(_02485_),
    .A2(_11833_),
    .B1(_11834_),
    .B2(_11835_),
    .X(_03108_));
 sky130_fd_sc_hd__buf_1 _15476_ (.A(pcpi_rs1[18]),
    .X(_11836_));
 sky130_fd_sc_hd__o22a_2 _15477_ (.A1(_02484_),
    .A2(_11833_),
    .B1(_11836_),
    .B2(_11835_),
    .X(_03107_));
 sky130_fd_sc_hd__buf_1 _15478_ (.A(pcpi_rs1[17]),
    .X(_11837_));
 sky130_fd_sc_hd__buf_1 _15479_ (.A(_11837_),
    .X(_11838_));
 sky130_fd_sc_hd__o22a_2 _15480_ (.A1(_02483_),
    .A2(_11833_),
    .B1(_11838_),
    .B2(_11835_),
    .X(_03106_));
 sky130_fd_sc_hd__buf_1 _15481_ (.A(pcpi_rs1[16]),
    .X(_11839_));
 sky130_fd_sc_hd__o22a_2 _15482_ (.A1(_02482_),
    .A2(_11833_),
    .B1(_11839_),
    .B2(_11835_),
    .X(_03105_));
 sky130_fd_sc_hd__buf_1 _15483_ (.A(pcpi_rs1[15]),
    .X(_11840_));
 sky130_fd_sc_hd__o22a_2 _15484_ (.A1(_02481_),
    .A2(_11833_),
    .B1(_11840_),
    .B2(_11835_),
    .X(_03104_));
 sky130_fd_sc_hd__buf_1 _15485_ (.A(pcpi_rs1[14]),
    .X(_11841_));
 sky130_fd_sc_hd__o22a_2 _15486_ (.A1(_02480_),
    .A2(_11833_),
    .B1(_11841_),
    .B2(_11835_),
    .X(_03103_));
 sky130_fd_sc_hd__buf_1 _15487_ (.A(_11810_),
    .X(_11842_));
 sky130_fd_sc_hd__buf_1 _15488_ (.A(pcpi_rs1[13]),
    .X(_11843_));
 sky130_fd_sc_hd__buf_1 _15489_ (.A(_11814_),
    .X(_11844_));
 sky130_fd_sc_hd__o22a_2 _15490_ (.A1(_02479_),
    .A2(_11842_),
    .B1(_11843_),
    .B2(_11844_),
    .X(_03102_));
 sky130_fd_sc_hd__buf_1 _15491_ (.A(pcpi_rs1[12]),
    .X(_11845_));
 sky130_fd_sc_hd__o22a_2 _15492_ (.A1(_02478_),
    .A2(_11842_),
    .B1(_11845_),
    .B2(_11844_),
    .X(_03101_));
 sky130_fd_sc_hd__buf_1 _15493_ (.A(pcpi_rs1[11]),
    .X(_11846_));
 sky130_fd_sc_hd__o22a_2 _15494_ (.A1(_02477_),
    .A2(_11842_),
    .B1(_11846_),
    .B2(_11844_),
    .X(_03100_));
 sky130_fd_sc_hd__buf_1 _15495_ (.A(pcpi_rs1[10]),
    .X(_11847_));
 sky130_fd_sc_hd__o22a_2 _15496_ (.A1(_02476_),
    .A2(_11842_),
    .B1(_11847_),
    .B2(_11844_),
    .X(_03099_));
 sky130_fd_sc_hd__buf_1 _15497_ (.A(pcpi_rs1[9]),
    .X(_11848_));
 sky130_fd_sc_hd__buf_1 _15498_ (.A(_11848_),
    .X(_11849_));
 sky130_fd_sc_hd__o22a_2 _15499_ (.A1(_02506_),
    .A2(_11842_),
    .B1(_11849_),
    .B2(_11844_),
    .X(_03098_));
 sky130_fd_sc_hd__buf_1 _15500_ (.A(pcpi_rs1[8]),
    .X(_11850_));
 sky130_fd_sc_hd__o22a_2 _15501_ (.A1(_02505_),
    .A2(_11842_),
    .B1(_11850_),
    .B2(_11844_),
    .X(_03097_));
 sky130_fd_sc_hd__buf_1 _15502_ (.A(_11809_),
    .X(_11851_));
 sky130_fd_sc_hd__buf_1 _15503_ (.A(pcpi_rs1[7]),
    .X(_11852_));
 sky130_fd_sc_hd__buf_1 _15504_ (.A(_11852_),
    .X(_11853_));
 sky130_fd_sc_hd__buf_1 _15505_ (.A(_11813_),
    .X(_11854_));
 sky130_fd_sc_hd__o22a_2 _15506_ (.A1(_02504_),
    .A2(_11851_),
    .B1(_11853_),
    .B2(_11854_),
    .X(_03096_));
 sky130_fd_sc_hd__buf_1 _15507_ (.A(pcpi_rs1[6]),
    .X(_11855_));
 sky130_fd_sc_hd__buf_1 _15508_ (.A(_11855_),
    .X(_11856_));
 sky130_fd_sc_hd__o22a_2 _15509_ (.A1(_02503_),
    .A2(_11851_),
    .B1(_11856_),
    .B2(_11854_),
    .X(_03095_));
 sky130_fd_sc_hd__buf_1 _15510_ (.A(pcpi_rs1[5]),
    .X(_11857_));
 sky130_fd_sc_hd__o22a_2 _15511_ (.A1(_02502_),
    .A2(_11851_),
    .B1(_11857_),
    .B2(_11854_),
    .X(_03094_));
 sky130_fd_sc_hd__buf_1 _15512_ (.A(pcpi_rs1[4]),
    .X(_11858_));
 sky130_fd_sc_hd__o22a_2 _15513_ (.A1(_02501_),
    .A2(_11851_),
    .B1(_11858_),
    .B2(_11854_),
    .X(_03093_));
 sky130_fd_sc_hd__buf_1 _15514_ (.A(pcpi_rs1[3]),
    .X(_11859_));
 sky130_fd_sc_hd__o22a_2 _15515_ (.A1(_02500_),
    .A2(_11851_),
    .B1(_11859_),
    .B2(_11854_),
    .X(_03092_));
 sky130_fd_sc_hd__buf_1 _15516_ (.A(pcpi_rs1[2]),
    .X(_11860_));
 sky130_fd_sc_hd__o22a_2 _15517_ (.A1(_02497_),
    .A2(_11851_),
    .B1(_11860_),
    .B2(_11854_),
    .X(_03091_));
 sky130_fd_sc_hd__buf_1 _15518_ (.A(pcpi_rs1[1]),
    .X(_11861_));
 sky130_fd_sc_hd__buf_1 _15519_ (.A(_11861_),
    .X(_11862_));
 sky130_fd_sc_hd__o22a_2 _15520_ (.A1(_02486_),
    .A2(_11810_),
    .B1(_11862_),
    .B2(_11814_),
    .X(_03090_));
 sky130_fd_sc_hd__buf_1 _15521_ (.A(pcpi_rs1[0]),
    .X(_11863_));
 sky130_fd_sc_hd__o22a_2 _15522_ (.A1(_02475_),
    .A2(_11810_),
    .B1(_11863_),
    .B2(_11814_),
    .X(_03089_));
 sky130_fd_sc_hd__buf_1 _15523_ (.A(_10710_),
    .X(_11864_));
 sky130_fd_sc_hd__a22o_2 _15524_ (.A1(mem_addr[31]),
    .A2(_10712_),
    .B1(mem_la_addr[31]),
    .B2(_11864_),
    .X(_03088_));
 sky130_fd_sc_hd__a22o_2 _15525_ (.A1(mem_addr[30]),
    .A2(_10712_),
    .B1(mem_la_addr[30]),
    .B2(_11864_),
    .X(_03087_));
 sky130_fd_sc_hd__a22o_2 _15526_ (.A1(mem_addr[29]),
    .A2(_10712_),
    .B1(mem_la_addr[29]),
    .B2(_11864_),
    .X(_03086_));
 sky130_fd_sc_hd__a22o_2 _15527_ (.A1(mem_addr[28]),
    .A2(_10712_),
    .B1(mem_la_addr[28]),
    .B2(_11864_),
    .X(_03085_));
 sky130_fd_sc_hd__a22o_2 _15528_ (.A1(mem_addr[27]),
    .A2(_10712_),
    .B1(mem_la_addr[27]),
    .B2(_11864_),
    .X(_03084_));
 sky130_fd_sc_hd__buf_1 _15529_ (.A(_10711_),
    .X(_11865_));
 sky130_fd_sc_hd__a22o_2 _15530_ (.A1(mem_addr[26]),
    .A2(_11865_),
    .B1(mem_la_addr[26]),
    .B2(_11864_),
    .X(_03083_));
 sky130_fd_sc_hd__buf_1 _15531_ (.A(_10710_),
    .X(_11866_));
 sky130_fd_sc_hd__a22o_2 _15532_ (.A1(mem_addr[25]),
    .A2(_11865_),
    .B1(mem_la_addr[25]),
    .B2(_11866_),
    .X(_03082_));
 sky130_fd_sc_hd__a22o_2 _15533_ (.A1(mem_addr[24]),
    .A2(_11865_),
    .B1(mem_la_addr[24]),
    .B2(_11866_),
    .X(_03081_));
 sky130_fd_sc_hd__a22o_2 _15534_ (.A1(mem_addr[23]),
    .A2(_11865_),
    .B1(mem_la_addr[23]),
    .B2(_11866_),
    .X(_03080_));
 sky130_fd_sc_hd__a22o_2 _15535_ (.A1(mem_addr[22]),
    .A2(_11865_),
    .B1(mem_la_addr[22]),
    .B2(_11866_),
    .X(_03079_));
 sky130_fd_sc_hd__a22o_2 _15536_ (.A1(mem_addr[21]),
    .A2(_11865_),
    .B1(mem_la_addr[21]),
    .B2(_11866_),
    .X(_03078_));
 sky130_fd_sc_hd__buf_1 _15537_ (.A(_10711_),
    .X(_11867_));
 sky130_fd_sc_hd__a22o_2 _15538_ (.A1(mem_addr[20]),
    .A2(_11867_),
    .B1(mem_la_addr[20]),
    .B2(_11866_),
    .X(_03077_));
 sky130_fd_sc_hd__buf_1 _15539_ (.A(_10710_),
    .X(_11868_));
 sky130_fd_sc_hd__a22o_2 _15540_ (.A1(mem_addr[19]),
    .A2(_11867_),
    .B1(mem_la_addr[19]),
    .B2(_11868_),
    .X(_03076_));
 sky130_fd_sc_hd__a22o_2 _15541_ (.A1(mem_addr[18]),
    .A2(_11867_),
    .B1(mem_la_addr[18]),
    .B2(_11868_),
    .X(_03075_));
 sky130_fd_sc_hd__a22o_2 _15542_ (.A1(mem_addr[17]),
    .A2(_11867_),
    .B1(mem_la_addr[17]),
    .B2(_11868_),
    .X(_03074_));
 sky130_fd_sc_hd__a22o_2 _15543_ (.A1(mem_addr[16]),
    .A2(_11867_),
    .B1(mem_la_addr[16]),
    .B2(_11868_),
    .X(_03073_));
 sky130_fd_sc_hd__a22o_2 _15544_ (.A1(mem_addr[15]),
    .A2(_11867_),
    .B1(mem_la_addr[15]),
    .B2(_11868_),
    .X(_03072_));
 sky130_fd_sc_hd__buf_1 _15545_ (.A(_10711_),
    .X(_11869_));
 sky130_fd_sc_hd__a22o_2 _15546_ (.A1(mem_addr[14]),
    .A2(_11869_),
    .B1(mem_la_addr[14]),
    .B2(_11868_),
    .X(_03071_));
 sky130_fd_sc_hd__buf_1 _15547_ (.A(_10710_),
    .X(_11870_));
 sky130_fd_sc_hd__a22o_2 _15548_ (.A1(mem_addr[13]),
    .A2(_11869_),
    .B1(mem_la_addr[13]),
    .B2(_11870_),
    .X(_03070_));
 sky130_fd_sc_hd__a22o_2 _15549_ (.A1(mem_addr[12]),
    .A2(_11869_),
    .B1(mem_la_addr[12]),
    .B2(_11870_),
    .X(_03069_));
 sky130_fd_sc_hd__a22o_2 _15550_ (.A1(mem_addr[11]),
    .A2(_11869_),
    .B1(mem_la_addr[11]),
    .B2(_11870_),
    .X(_03068_));
 sky130_fd_sc_hd__a22o_2 _15551_ (.A1(mem_addr[10]),
    .A2(_11869_),
    .B1(mem_la_addr[10]),
    .B2(_11870_),
    .X(_03067_));
 sky130_fd_sc_hd__a22o_2 _15552_ (.A1(mem_addr[9]),
    .A2(_11869_),
    .B1(mem_la_addr[9]),
    .B2(_11870_),
    .X(_03066_));
 sky130_fd_sc_hd__buf_1 _15553_ (.A(_10711_),
    .X(_11871_));
 sky130_fd_sc_hd__a22o_2 _15554_ (.A1(mem_addr[8]),
    .A2(_11871_),
    .B1(mem_la_addr[8]),
    .B2(_11870_),
    .X(_03065_));
 sky130_fd_sc_hd__buf_1 _15555_ (.A(_10710_),
    .X(_11872_));
 sky130_fd_sc_hd__a22o_2 _15556_ (.A1(mem_addr[7]),
    .A2(_11871_),
    .B1(mem_la_addr[7]),
    .B2(_11872_),
    .X(_03064_));
 sky130_fd_sc_hd__a22o_2 _15557_ (.A1(mem_addr[6]),
    .A2(_11871_),
    .B1(mem_la_addr[6]),
    .B2(_11872_),
    .X(_03063_));
 sky130_fd_sc_hd__a22o_2 _15558_ (.A1(mem_addr[5]),
    .A2(_11871_),
    .B1(mem_la_addr[5]),
    .B2(_11872_),
    .X(_03062_));
 sky130_fd_sc_hd__a22o_2 _15559_ (.A1(mem_addr[4]),
    .A2(_11871_),
    .B1(mem_la_addr[4]),
    .B2(_11872_),
    .X(_03061_));
 sky130_fd_sc_hd__a22o_2 _15560_ (.A1(mem_addr[3]),
    .A2(_11871_),
    .B1(mem_la_addr[3]),
    .B2(_11872_),
    .X(_03060_));
 sky130_fd_sc_hd__a22o_2 _15561_ (.A1(mem_addr[2]),
    .A2(_10711_),
    .B1(mem_la_addr[2]),
    .B2(_11872_),
    .X(_03059_));
 sky130_fd_sc_hd__buf_1 _15562_ (.A(\pcpi_mul.rs1[31] ),
    .X(_11873_));
 sky130_fd_sc_hd__buf_1 _15563_ (.A(_11873_),
    .X(_11874_));
 sky130_fd_sc_hd__buf_1 _15564_ (.A(_11874_),
    .X(_11875_));
 sky130_fd_sc_hd__a22o_2 _15565_ (.A1(_11812_),
    .A2(_10592_),
    .B1(_11875_),
    .B2(_11565_),
    .X(_03058_));
 sky130_fd_sc_hd__buf_1 _15566_ (.A(\pcpi_mul.rs1[30] ),
    .X(_11876_));
 sky130_fd_sc_hd__buf_1 _15567_ (.A(_11876_),
    .X(_11877_));
 sky130_fd_sc_hd__buf_1 _15568_ (.A(_11877_),
    .X(_11878_));
 sky130_fd_sc_hd__buf_1 _15569_ (.A(_11878_),
    .X(_11879_));
 sky130_fd_sc_hd__a22o_2 _15570_ (.A1(_11879_),
    .A2(_11639_),
    .B1(_11816_),
    .B2(_11645_),
    .X(_03057_));
 sky130_fd_sc_hd__buf_1 _15571_ (.A(\pcpi_mul.rs1[29] ),
    .X(_11880_));
 sky130_fd_sc_hd__buf_1 _15572_ (.A(_11880_),
    .X(_11881_));
 sky130_fd_sc_hd__a22o_2 _15573_ (.A1(_11881_),
    .A2(_11639_),
    .B1(_11817_),
    .B2(_11645_),
    .X(_03056_));
 sky130_fd_sc_hd__buf_1 _15574_ (.A(\pcpi_mul.rs1[28] ),
    .X(_11882_));
 sky130_fd_sc_hd__buf_1 _15575_ (.A(_11882_),
    .X(_11883_));
 sky130_fd_sc_hd__a22o_2 _15576_ (.A1(_11883_),
    .A2(_11639_),
    .B1(_11818_),
    .B2(_11645_),
    .X(_03055_));
 sky130_fd_sc_hd__buf_1 _15577_ (.A(\pcpi_mul.rs1[27] ),
    .X(_11884_));
 sky130_fd_sc_hd__buf_1 _15578_ (.A(_11884_),
    .X(_11885_));
 sky130_fd_sc_hd__buf_1 _15579_ (.A(_11885_),
    .X(_11886_));
 sky130_fd_sc_hd__buf_1 _15580_ (.A(_11595_),
    .X(_11887_));
 sky130_fd_sc_hd__a22o_2 _15581_ (.A1(_11886_),
    .A2(_11887_),
    .B1(_11820_),
    .B2(_11645_),
    .X(_03054_));
 sky130_fd_sc_hd__buf_1 _15582_ (.A(\pcpi_mul.rs1[26] ),
    .X(_11888_));
 sky130_fd_sc_hd__buf_1 _15583_ (.A(_11888_),
    .X(_11889_));
 sky130_fd_sc_hd__buf_1 _15584_ (.A(_11889_),
    .X(_11890_));
 sky130_fd_sc_hd__buf_1 _15585_ (.A(_10591_),
    .X(_11891_));
 sky130_fd_sc_hd__a22o_2 _15586_ (.A1(_11890_),
    .A2(_11887_),
    .B1(_11822_),
    .B2(_11891_),
    .X(_03053_));
 sky130_fd_sc_hd__buf_1 _15587_ (.A(\pcpi_mul.rs1[25] ),
    .X(_11892_));
 sky130_fd_sc_hd__buf_1 _15588_ (.A(_11892_),
    .X(_11893_));
 sky130_fd_sc_hd__buf_1 _15589_ (.A(_11893_),
    .X(_11894_));
 sky130_fd_sc_hd__a22o_2 _15590_ (.A1(_11894_),
    .A2(_11887_),
    .B1(_11825_),
    .B2(_11891_),
    .X(_03052_));
 sky130_fd_sc_hd__buf_1 _15591_ (.A(\pcpi_mul.rs1[24] ),
    .X(_11895_));
 sky130_fd_sc_hd__buf_1 _15592_ (.A(_11895_),
    .X(_11896_));
 sky130_fd_sc_hd__a22o_2 _15593_ (.A1(_11896_),
    .A2(_11887_),
    .B1(_11828_),
    .B2(_11891_),
    .X(_03051_));
 sky130_fd_sc_hd__buf_1 _15594_ (.A(\pcpi_mul.rs1[23] ),
    .X(_11897_));
 sky130_fd_sc_hd__buf_1 _15595_ (.A(_11897_),
    .X(_11898_));
 sky130_fd_sc_hd__a22o_2 _15596_ (.A1(_11898_),
    .A2(_11887_),
    .B1(_11829_),
    .B2(_11891_),
    .X(_03050_));
 sky130_fd_sc_hd__buf_1 _15597_ (.A(\pcpi_mul.rs1[22] ),
    .X(_11899_));
 sky130_fd_sc_hd__buf_1 _15598_ (.A(_11899_),
    .X(_11900_));
 sky130_fd_sc_hd__buf_1 _15599_ (.A(_11900_),
    .X(_11901_));
 sky130_fd_sc_hd__a22o_2 _15600_ (.A1(_11901_),
    .A2(_11887_),
    .B1(_11830_),
    .B2(_11891_),
    .X(_03049_));
 sky130_fd_sc_hd__buf_1 _15601_ (.A(\pcpi_mul.rs1[21] ),
    .X(_11902_));
 sky130_fd_sc_hd__buf_1 _15602_ (.A(_11902_),
    .X(_11903_));
 sky130_fd_sc_hd__buf_1 _15603_ (.A(_11595_),
    .X(_11904_));
 sky130_fd_sc_hd__a22o_2 _15604_ (.A1(_11903_),
    .A2(_11904_),
    .B1(_11831_),
    .B2(_11891_),
    .X(_03048_));
 sky130_fd_sc_hd__buf_1 _15605_ (.A(\pcpi_mul.rs1[20] ),
    .X(_11905_));
 sky130_fd_sc_hd__buf_1 _15606_ (.A(_11905_),
    .X(_11906_));
 sky130_fd_sc_hd__buf_1 _15607_ (.A(_10591_),
    .X(_11907_));
 sky130_fd_sc_hd__a22o_2 _15608_ (.A1(_11906_),
    .A2(_11904_),
    .B1(_11832_),
    .B2(_11907_),
    .X(_03047_));
 sky130_fd_sc_hd__buf_1 _15609_ (.A(\pcpi_mul.rs1[19] ),
    .X(_11908_));
 sky130_fd_sc_hd__buf_1 _15610_ (.A(_11908_),
    .X(_11909_));
 sky130_fd_sc_hd__a22o_2 _15611_ (.A1(_11909_),
    .A2(_11904_),
    .B1(_11834_),
    .B2(_11907_),
    .X(_03046_));
 sky130_fd_sc_hd__buf_1 _15612_ (.A(\pcpi_mul.rs1[18] ),
    .X(_11910_));
 sky130_fd_sc_hd__buf_1 _15613_ (.A(_11910_),
    .X(_11911_));
 sky130_fd_sc_hd__a22o_2 _15614_ (.A1(_11911_),
    .A2(_11904_),
    .B1(_11836_),
    .B2(_11907_),
    .X(_03045_));
 sky130_fd_sc_hd__buf_1 _15615_ (.A(\pcpi_mul.rs1[17] ),
    .X(_11912_));
 sky130_fd_sc_hd__buf_1 _15616_ (.A(_11912_),
    .X(_11913_));
 sky130_fd_sc_hd__a22o_2 _15617_ (.A1(_11913_),
    .A2(_11904_),
    .B1(_11838_),
    .B2(_11907_),
    .X(_03044_));
 sky130_fd_sc_hd__buf_1 _15618_ (.A(\pcpi_mul.rs1[16] ),
    .X(_11914_));
 sky130_fd_sc_hd__buf_1 _15619_ (.A(_11914_),
    .X(_11915_));
 sky130_fd_sc_hd__a22o_2 _15620_ (.A1(_11915_),
    .A2(_11904_),
    .B1(_11839_),
    .B2(_11907_),
    .X(_03043_));
 sky130_fd_sc_hd__buf_1 _15621_ (.A(\pcpi_mul.rs1[15] ),
    .X(_11916_));
 sky130_fd_sc_hd__buf_1 _15622_ (.A(_11916_),
    .X(_11917_));
 sky130_fd_sc_hd__buf_1 _15623_ (.A(_10578_),
    .X(_11918_));
 sky130_fd_sc_hd__a22o_2 _15624_ (.A1(_11917_),
    .A2(_11918_),
    .B1(_11840_),
    .B2(_11907_),
    .X(_03042_));
 sky130_fd_sc_hd__buf_1 _15625_ (.A(\pcpi_mul.rs1[14] ),
    .X(_11919_));
 sky130_fd_sc_hd__buf_1 _15626_ (.A(_11919_),
    .X(_11920_));
 sky130_fd_sc_hd__buf_1 _15627_ (.A(_10591_),
    .X(_11921_));
 sky130_fd_sc_hd__a22o_2 _15628_ (.A1(_11920_),
    .A2(_11918_),
    .B1(_11841_),
    .B2(_11921_),
    .X(_03041_));
 sky130_fd_sc_hd__buf_1 _15629_ (.A(\pcpi_mul.rs1[13] ),
    .X(_11922_));
 sky130_fd_sc_hd__buf_1 _15630_ (.A(_11922_),
    .X(_11923_));
 sky130_fd_sc_hd__a22o_2 _15631_ (.A1(_11923_),
    .A2(_11918_),
    .B1(_11843_),
    .B2(_11921_),
    .X(_03040_));
 sky130_fd_sc_hd__buf_1 _15632_ (.A(\pcpi_mul.rs1[12] ),
    .X(_11924_));
 sky130_fd_sc_hd__buf_1 _15633_ (.A(_11924_),
    .X(_11925_));
 sky130_fd_sc_hd__a22o_2 _15634_ (.A1(_11925_),
    .A2(_11918_),
    .B1(_11845_),
    .B2(_11921_),
    .X(_03039_));
 sky130_fd_sc_hd__buf_1 _15635_ (.A(\pcpi_mul.rs1[11] ),
    .X(_11926_));
 sky130_fd_sc_hd__buf_1 _15636_ (.A(_11926_),
    .X(_11927_));
 sky130_fd_sc_hd__a22o_2 _15637_ (.A1(_11927_),
    .A2(_11918_),
    .B1(_11846_),
    .B2(_11921_),
    .X(_03038_));
 sky130_fd_sc_hd__buf_1 _15638_ (.A(\pcpi_mul.rs1[10] ),
    .X(_11928_));
 sky130_fd_sc_hd__buf_1 _15639_ (.A(_11928_),
    .X(_11929_));
 sky130_fd_sc_hd__a22o_2 _15640_ (.A1(_11929_),
    .A2(_11918_),
    .B1(_11847_),
    .B2(_11921_),
    .X(_03037_));
 sky130_fd_sc_hd__buf_1 _15641_ (.A(\pcpi_mul.rs1[9] ),
    .X(_11930_));
 sky130_fd_sc_hd__buf_1 _15642_ (.A(_11930_),
    .X(_11931_));
 sky130_fd_sc_hd__buf_1 _15643_ (.A(_10578_),
    .X(_11932_));
 sky130_fd_sc_hd__a22o_2 _15644_ (.A1(_11931_),
    .A2(_11932_),
    .B1(_11849_),
    .B2(_11921_),
    .X(_03036_));
 sky130_fd_sc_hd__buf_1 _15645_ (.A(\pcpi_mul.rs1[8] ),
    .X(_11933_));
 sky130_fd_sc_hd__buf_1 _15646_ (.A(_11933_),
    .X(_11934_));
 sky130_fd_sc_hd__buf_1 _15647_ (.A(_10591_),
    .X(_11935_));
 sky130_fd_sc_hd__a22o_2 _15648_ (.A1(_11934_),
    .A2(_11932_),
    .B1(_11850_),
    .B2(_11935_),
    .X(_03035_));
 sky130_fd_sc_hd__buf_1 _15649_ (.A(\pcpi_mul.rs1[7] ),
    .X(_11936_));
 sky130_fd_sc_hd__buf_1 _15650_ (.A(_11936_),
    .X(_11937_));
 sky130_fd_sc_hd__a22o_2 _15651_ (.A1(_11937_),
    .A2(_11932_),
    .B1(_11853_),
    .B2(_11935_),
    .X(_03034_));
 sky130_fd_sc_hd__buf_1 _15652_ (.A(\pcpi_mul.rs1[6] ),
    .X(_11938_));
 sky130_fd_sc_hd__buf_1 _15653_ (.A(_11938_),
    .X(_11939_));
 sky130_fd_sc_hd__buf_1 _15654_ (.A(_11939_),
    .X(_11940_));
 sky130_fd_sc_hd__a22o_2 _15655_ (.A1(_11940_),
    .A2(_11932_),
    .B1(_11856_),
    .B2(_11935_),
    .X(_03033_));
 sky130_fd_sc_hd__buf_1 _15656_ (.A(\pcpi_mul.rs1[5] ),
    .X(_11941_));
 sky130_fd_sc_hd__buf_1 _15657_ (.A(_11941_),
    .X(_11942_));
 sky130_fd_sc_hd__buf_1 _15658_ (.A(_11942_),
    .X(_11943_));
 sky130_fd_sc_hd__a22o_2 _15659_ (.A1(_11943_),
    .A2(_11932_),
    .B1(_11857_),
    .B2(_11935_),
    .X(_03032_));
 sky130_fd_sc_hd__buf_1 _15660_ (.A(\pcpi_mul.rs1[4] ),
    .X(_11944_));
 sky130_fd_sc_hd__buf_1 _15661_ (.A(_11944_),
    .X(_11945_));
 sky130_fd_sc_hd__buf_1 _15662_ (.A(_11945_),
    .X(_11946_));
 sky130_fd_sc_hd__a22o_2 _15663_ (.A1(_11946_),
    .A2(_11932_),
    .B1(_11858_),
    .B2(_11935_),
    .X(_03031_));
 sky130_fd_sc_hd__buf_1 _15664_ (.A(\pcpi_mul.rs1[3] ),
    .X(_11947_));
 sky130_fd_sc_hd__buf_1 _15665_ (.A(_11947_),
    .X(_11948_));
 sky130_fd_sc_hd__buf_1 _15666_ (.A(_11948_),
    .X(_11949_));
 sky130_fd_sc_hd__a22o_2 _15667_ (.A1(_11949_),
    .A2(_11564_),
    .B1(_11859_),
    .B2(_11935_),
    .X(_03030_));
 sky130_fd_sc_hd__buf_1 _15668_ (.A(\pcpi_mul.rs1[2] ),
    .X(_11950_));
 sky130_fd_sc_hd__buf_1 _15669_ (.A(_11950_),
    .X(_11951_));
 sky130_fd_sc_hd__buf_1 _15670_ (.A(_11951_),
    .X(_11952_));
 sky130_fd_sc_hd__a22o_2 _15671_ (.A1(_11952_),
    .A2(_11564_),
    .B1(_11860_),
    .B2(_10592_),
    .X(_03029_));
 sky130_fd_sc_hd__buf_1 _15672_ (.A(\pcpi_mul.rs1[1] ),
    .X(_11953_));
 sky130_fd_sc_hd__buf_1 _15673_ (.A(_11953_),
    .X(_11954_));
 sky130_fd_sc_hd__buf_1 _15674_ (.A(_11954_),
    .X(_11955_));
 sky130_fd_sc_hd__a22o_2 _15675_ (.A1(_11955_),
    .A2(_11564_),
    .B1(_11862_),
    .B2(_10592_),
    .X(_03028_));
 sky130_fd_sc_hd__buf_1 _15676_ (.A(\pcpi_mul.rs1[0] ),
    .X(_11956_));
 sky130_fd_sc_hd__buf_1 _15677_ (.A(_11956_),
    .X(_11957_));
 sky130_fd_sc_hd__a22o_2 _15678_ (.A1(_11957_),
    .A2(_11564_),
    .B1(_11863_),
    .B2(_10592_),
    .X(_03027_));
 sky130_fd_sc_hd__or2_2 _15679_ (.A(_11254_),
    .B(_11313_),
    .X(_11958_));
 sky130_fd_sc_hd__buf_1 _15680_ (.A(_11958_),
    .X(_11959_));
 sky130_fd_sc_hd__buf_1 _15681_ (.A(_11959_),
    .X(_11960_));
 sky130_vsdinv _15682_ (.A(_11958_),
    .Y(_11961_));
 sky130_fd_sc_hd__buf_1 _15683_ (.A(_11961_),
    .X(_11962_));
 sky130_fd_sc_hd__buf_1 _15684_ (.A(_11962_),
    .X(_11963_));
 sky130_fd_sc_hd__a22o_2 _15685_ (.A1(\cpuregs[5][31] ),
    .A2(_11960_),
    .B1(_11653_),
    .B2(_11963_),
    .X(_03026_));
 sky130_fd_sc_hd__a22o_2 _15686_ (.A1(\cpuregs[5][30] ),
    .A2(_11960_),
    .B1(_11657_),
    .B2(_11963_),
    .X(_03025_));
 sky130_fd_sc_hd__a22o_2 _15687_ (.A1(\cpuregs[5][29] ),
    .A2(_11960_),
    .B1(_11658_),
    .B2(_11963_),
    .X(_03024_));
 sky130_fd_sc_hd__a22o_2 _15688_ (.A1(\cpuregs[5][28] ),
    .A2(_11960_),
    .B1(_11659_),
    .B2(_11963_),
    .X(_03023_));
 sky130_fd_sc_hd__a22o_2 _15689_ (.A1(\cpuregs[5][27] ),
    .A2(_11960_),
    .B1(_11660_),
    .B2(_11963_),
    .X(_03022_));
 sky130_fd_sc_hd__a22o_2 _15690_ (.A1(\cpuregs[5][26] ),
    .A2(_11960_),
    .B1(_11661_),
    .B2(_11963_),
    .X(_03021_));
 sky130_fd_sc_hd__buf_1 _15691_ (.A(_11959_),
    .X(_11964_));
 sky130_fd_sc_hd__buf_1 _15692_ (.A(_11962_),
    .X(_11965_));
 sky130_fd_sc_hd__a22o_2 _15693_ (.A1(\cpuregs[5][25] ),
    .A2(_11964_),
    .B1(_11663_),
    .B2(_11965_),
    .X(_03020_));
 sky130_fd_sc_hd__a22o_2 _15694_ (.A1(\cpuregs[5][24] ),
    .A2(_11964_),
    .B1(_11665_),
    .B2(_11965_),
    .X(_03019_));
 sky130_fd_sc_hd__a22o_2 _15695_ (.A1(\cpuregs[5][23] ),
    .A2(_11964_),
    .B1(_11666_),
    .B2(_11965_),
    .X(_03018_));
 sky130_fd_sc_hd__a22o_2 _15696_ (.A1(\cpuregs[5][22] ),
    .A2(_11964_),
    .B1(_11667_),
    .B2(_11965_),
    .X(_03017_));
 sky130_fd_sc_hd__a22o_2 _15697_ (.A1(\cpuregs[5][21] ),
    .A2(_11964_),
    .B1(_11668_),
    .B2(_11965_),
    .X(_03016_));
 sky130_fd_sc_hd__a22o_2 _15698_ (.A1(\cpuregs[5][20] ),
    .A2(_11964_),
    .B1(_11669_),
    .B2(_11965_),
    .X(_03015_));
 sky130_fd_sc_hd__buf_1 _15699_ (.A(_11959_),
    .X(_11966_));
 sky130_fd_sc_hd__buf_1 _15700_ (.A(_11962_),
    .X(_11967_));
 sky130_fd_sc_hd__a22o_2 _15701_ (.A1(\cpuregs[5][19] ),
    .A2(_11966_),
    .B1(_11671_),
    .B2(_11967_),
    .X(_03014_));
 sky130_fd_sc_hd__a22o_2 _15702_ (.A1(\cpuregs[5][18] ),
    .A2(_11966_),
    .B1(_11673_),
    .B2(_11967_),
    .X(_03013_));
 sky130_fd_sc_hd__a22o_2 _15703_ (.A1(\cpuregs[5][17] ),
    .A2(_11966_),
    .B1(_11674_),
    .B2(_11967_),
    .X(_03012_));
 sky130_fd_sc_hd__a22o_2 _15704_ (.A1(\cpuregs[5][16] ),
    .A2(_11966_),
    .B1(_11675_),
    .B2(_11967_),
    .X(_03011_));
 sky130_fd_sc_hd__a22o_2 _15705_ (.A1(\cpuregs[5][15] ),
    .A2(_11966_),
    .B1(_11676_),
    .B2(_11967_),
    .X(_03010_));
 sky130_fd_sc_hd__a22o_2 _15706_ (.A1(\cpuregs[5][14] ),
    .A2(_11966_),
    .B1(_11677_),
    .B2(_11967_),
    .X(_03009_));
 sky130_fd_sc_hd__buf_1 _15707_ (.A(_11959_),
    .X(_11968_));
 sky130_fd_sc_hd__buf_1 _15708_ (.A(_11962_),
    .X(_11969_));
 sky130_fd_sc_hd__a22o_2 _15709_ (.A1(\cpuregs[5][13] ),
    .A2(_11968_),
    .B1(_11679_),
    .B2(_11969_),
    .X(_03008_));
 sky130_fd_sc_hd__a22o_2 _15710_ (.A1(\cpuregs[5][12] ),
    .A2(_11968_),
    .B1(_11681_),
    .B2(_11969_),
    .X(_03007_));
 sky130_fd_sc_hd__a22o_2 _15711_ (.A1(\cpuregs[5][11] ),
    .A2(_11968_),
    .B1(_11682_),
    .B2(_11969_),
    .X(_03006_));
 sky130_fd_sc_hd__a22o_2 _15712_ (.A1(\cpuregs[5][10] ),
    .A2(_11968_),
    .B1(_11683_),
    .B2(_11969_),
    .X(_03005_));
 sky130_fd_sc_hd__a22o_2 _15713_ (.A1(\cpuregs[5][9] ),
    .A2(_11968_),
    .B1(_11684_),
    .B2(_11969_),
    .X(_03004_));
 sky130_fd_sc_hd__a22o_2 _15714_ (.A1(\cpuregs[5][8] ),
    .A2(_11968_),
    .B1(_11685_),
    .B2(_11969_),
    .X(_03003_));
 sky130_fd_sc_hd__buf_1 _15715_ (.A(_11958_),
    .X(_11970_));
 sky130_fd_sc_hd__buf_1 _15716_ (.A(_11961_),
    .X(_11971_));
 sky130_fd_sc_hd__a22o_2 _15717_ (.A1(\cpuregs[5][7] ),
    .A2(_11970_),
    .B1(_11687_),
    .B2(_11971_),
    .X(_03002_));
 sky130_fd_sc_hd__a22o_2 _15718_ (.A1(\cpuregs[5][6] ),
    .A2(_11970_),
    .B1(_11689_),
    .B2(_11971_),
    .X(_03001_));
 sky130_fd_sc_hd__a22o_2 _15719_ (.A1(\cpuregs[5][5] ),
    .A2(_11970_),
    .B1(_11690_),
    .B2(_11971_),
    .X(_03000_));
 sky130_fd_sc_hd__a22o_2 _15720_ (.A1(\cpuregs[5][4] ),
    .A2(_11970_),
    .B1(_11691_),
    .B2(_11971_),
    .X(_02999_));
 sky130_fd_sc_hd__a22o_2 _15721_ (.A1(\cpuregs[5][3] ),
    .A2(_11970_),
    .B1(_11692_),
    .B2(_11971_),
    .X(_02998_));
 sky130_fd_sc_hd__a22o_2 _15722_ (.A1(\cpuregs[5][2] ),
    .A2(_11970_),
    .B1(_11693_),
    .B2(_11971_),
    .X(_02997_));
 sky130_fd_sc_hd__a22o_2 _15723_ (.A1(\cpuregs[5][1] ),
    .A2(_11959_),
    .B1(_11694_),
    .B2(_11962_),
    .X(_02996_));
 sky130_fd_sc_hd__a22o_2 _15724_ (.A1(\cpuregs[5][0] ),
    .A2(_11959_),
    .B1(_11695_),
    .B2(_11962_),
    .X(_02995_));
 sky130_fd_sc_hd__or2_2 _15725_ (.A(_11258_),
    .B(_11262_),
    .X(_11972_));
 sky130_fd_sc_hd__buf_1 _15726_ (.A(_11972_),
    .X(_11973_));
 sky130_fd_sc_hd__buf_1 _15727_ (.A(_11973_),
    .X(_11974_));
 sky130_vsdinv _15728_ (.A(_11972_),
    .Y(_11975_));
 sky130_fd_sc_hd__buf_1 _15729_ (.A(_11975_),
    .X(_11976_));
 sky130_fd_sc_hd__buf_1 _15730_ (.A(_11976_),
    .X(_11977_));
 sky130_fd_sc_hd__a22o_2 _15731_ (.A1(\cpuregs[2][31] ),
    .A2(_11974_),
    .B1(_11653_),
    .B2(_11977_),
    .X(_02994_));
 sky130_fd_sc_hd__a22o_2 _15732_ (.A1(\cpuregs[2][30] ),
    .A2(_11974_),
    .B1(_11657_),
    .B2(_11977_),
    .X(_02993_));
 sky130_fd_sc_hd__a22o_2 _15733_ (.A1(\cpuregs[2][29] ),
    .A2(_11974_),
    .B1(_11658_),
    .B2(_11977_),
    .X(_02992_));
 sky130_fd_sc_hd__a22o_2 _15734_ (.A1(\cpuregs[2][28] ),
    .A2(_11974_),
    .B1(_11659_),
    .B2(_11977_),
    .X(_02991_));
 sky130_fd_sc_hd__a22o_2 _15735_ (.A1(\cpuregs[2][27] ),
    .A2(_11974_),
    .B1(_11660_),
    .B2(_11977_),
    .X(_02990_));
 sky130_fd_sc_hd__a22o_2 _15736_ (.A1(\cpuregs[2][26] ),
    .A2(_11974_),
    .B1(_11661_),
    .B2(_11977_),
    .X(_02989_));
 sky130_fd_sc_hd__buf_1 _15737_ (.A(_11973_),
    .X(_11978_));
 sky130_fd_sc_hd__buf_1 _15738_ (.A(_11976_),
    .X(_11979_));
 sky130_fd_sc_hd__a22o_2 _15739_ (.A1(\cpuregs[2][25] ),
    .A2(_11978_),
    .B1(_11663_),
    .B2(_11979_),
    .X(_02988_));
 sky130_fd_sc_hd__a22o_2 _15740_ (.A1(\cpuregs[2][24] ),
    .A2(_11978_),
    .B1(_11665_),
    .B2(_11979_),
    .X(_02987_));
 sky130_fd_sc_hd__a22o_2 _15741_ (.A1(\cpuregs[2][23] ),
    .A2(_11978_),
    .B1(_11666_),
    .B2(_11979_),
    .X(_02986_));
 sky130_fd_sc_hd__a22o_2 _15742_ (.A1(\cpuregs[2][22] ),
    .A2(_11978_),
    .B1(_11667_),
    .B2(_11979_),
    .X(_02985_));
 sky130_fd_sc_hd__a22o_2 _15743_ (.A1(\cpuregs[2][21] ),
    .A2(_11978_),
    .B1(_11668_),
    .B2(_11979_),
    .X(_02984_));
 sky130_fd_sc_hd__a22o_2 _15744_ (.A1(\cpuregs[2][20] ),
    .A2(_11978_),
    .B1(_11669_),
    .B2(_11979_),
    .X(_02983_));
 sky130_fd_sc_hd__buf_1 _15745_ (.A(_11973_),
    .X(_11980_));
 sky130_fd_sc_hd__buf_1 _15746_ (.A(_11976_),
    .X(_11981_));
 sky130_fd_sc_hd__a22o_2 _15747_ (.A1(\cpuregs[2][19] ),
    .A2(_11980_),
    .B1(_11671_),
    .B2(_11981_),
    .X(_02982_));
 sky130_fd_sc_hd__a22o_2 _15748_ (.A1(\cpuregs[2][18] ),
    .A2(_11980_),
    .B1(_11673_),
    .B2(_11981_),
    .X(_02981_));
 sky130_fd_sc_hd__a22o_2 _15749_ (.A1(\cpuregs[2][17] ),
    .A2(_11980_),
    .B1(_11674_),
    .B2(_11981_),
    .X(_02980_));
 sky130_fd_sc_hd__a22o_2 _15750_ (.A1(\cpuregs[2][16] ),
    .A2(_11980_),
    .B1(_11675_),
    .B2(_11981_),
    .X(_02979_));
 sky130_fd_sc_hd__a22o_2 _15751_ (.A1(\cpuregs[2][15] ),
    .A2(_11980_),
    .B1(_11676_),
    .B2(_11981_),
    .X(_02978_));
 sky130_fd_sc_hd__a22o_2 _15752_ (.A1(\cpuregs[2][14] ),
    .A2(_11980_),
    .B1(_11677_),
    .B2(_11981_),
    .X(_02977_));
 sky130_fd_sc_hd__buf_1 _15753_ (.A(_11973_),
    .X(_11982_));
 sky130_fd_sc_hd__buf_1 _15754_ (.A(_11976_),
    .X(_11983_));
 sky130_fd_sc_hd__a22o_2 _15755_ (.A1(\cpuregs[2][13] ),
    .A2(_11982_),
    .B1(_11679_),
    .B2(_11983_),
    .X(_02976_));
 sky130_fd_sc_hd__a22o_2 _15756_ (.A1(\cpuregs[2][12] ),
    .A2(_11982_),
    .B1(_11681_),
    .B2(_11983_),
    .X(_02975_));
 sky130_fd_sc_hd__a22o_2 _15757_ (.A1(\cpuregs[2][11] ),
    .A2(_11982_),
    .B1(_11682_),
    .B2(_11983_),
    .X(_02974_));
 sky130_fd_sc_hd__a22o_2 _15758_ (.A1(\cpuregs[2][10] ),
    .A2(_11982_),
    .B1(_11683_),
    .B2(_11983_),
    .X(_02973_));
 sky130_fd_sc_hd__a22o_2 _15759_ (.A1(\cpuregs[2][9] ),
    .A2(_11982_),
    .B1(_11684_),
    .B2(_11983_),
    .X(_02972_));
 sky130_fd_sc_hd__a22o_2 _15760_ (.A1(\cpuregs[2][8] ),
    .A2(_11982_),
    .B1(_11685_),
    .B2(_11983_),
    .X(_02971_));
 sky130_fd_sc_hd__buf_1 _15761_ (.A(_11972_),
    .X(_11984_));
 sky130_fd_sc_hd__buf_1 _15762_ (.A(_11975_),
    .X(_11985_));
 sky130_fd_sc_hd__a22o_2 _15763_ (.A1(\cpuregs[2][7] ),
    .A2(_11984_),
    .B1(_11687_),
    .B2(_11985_),
    .X(_02970_));
 sky130_fd_sc_hd__a22o_2 _15764_ (.A1(\cpuregs[2][6] ),
    .A2(_11984_),
    .B1(_11689_),
    .B2(_11985_),
    .X(_02969_));
 sky130_fd_sc_hd__a22o_2 _15765_ (.A1(\cpuregs[2][5] ),
    .A2(_11984_),
    .B1(_11690_),
    .B2(_11985_),
    .X(_02968_));
 sky130_fd_sc_hd__a22o_2 _15766_ (.A1(\cpuregs[2][4] ),
    .A2(_11984_),
    .B1(_11691_),
    .B2(_11985_),
    .X(_02967_));
 sky130_fd_sc_hd__a22o_2 _15767_ (.A1(\cpuregs[2][3] ),
    .A2(_11984_),
    .B1(_11692_),
    .B2(_11985_),
    .X(_02966_));
 sky130_fd_sc_hd__a22o_2 _15768_ (.A1(\cpuregs[2][2] ),
    .A2(_11984_),
    .B1(_11693_),
    .B2(_11985_),
    .X(_02965_));
 sky130_fd_sc_hd__a22o_2 _15769_ (.A1(\cpuregs[2][1] ),
    .A2(_11973_),
    .B1(_11694_),
    .B2(_11976_),
    .X(_02964_));
 sky130_fd_sc_hd__a22o_2 _15770_ (.A1(\cpuregs[2][0] ),
    .A2(_11973_),
    .B1(_11695_),
    .B2(_11976_),
    .X(_02963_));
 sky130_fd_sc_hd__buf_1 _15771_ (.A(_10447_),
    .X(_11986_));
 sky130_fd_sc_hd__buf_1 _15772_ (.A(_11986_),
    .X(mem_xfer));
 sky130_fd_sc_hd__buf_1 _15773_ (.A(_10445_),
    .X(_11987_));
 sky130_fd_sc_hd__buf_1 _15774_ (.A(_11987_),
    .X(_11988_));
 sky130_fd_sc_hd__a22o_2 _15775_ (.A1(_10742_),
    .A2(_11988_),
    .B1(mem_rdata[31]),
    .B2(mem_xfer),
    .X(_02962_));
 sky130_fd_sc_hd__a22o_2 _15776_ (.A1(\mem_rdata_q[30] ),
    .A2(_11988_),
    .B1(mem_rdata[30]),
    .B2(mem_xfer),
    .X(_02961_));
 sky130_fd_sc_hd__a22o_2 _15777_ (.A1(_10740_),
    .A2(_11988_),
    .B1(mem_rdata[29]),
    .B2(mem_xfer),
    .X(_02960_));
 sky130_fd_sc_hd__a22o_2 _15778_ (.A1(_11729_),
    .A2(_11988_),
    .B1(mem_rdata[28]),
    .B2(mem_xfer),
    .X(_02959_));
 sky130_fd_sc_hd__buf_1 _15779_ (.A(_11986_),
    .X(_11989_));
 sky130_fd_sc_hd__a22o_2 _15780_ (.A1(_11722_),
    .A2(_11988_),
    .B1(mem_rdata[27]),
    .B2(_11989_),
    .X(_02958_));
 sky130_fd_sc_hd__a22o_2 _15781_ (.A1(_11730_),
    .A2(_11988_),
    .B1(mem_rdata[26]),
    .B2(_11989_),
    .X(_02957_));
 sky130_fd_sc_hd__buf_1 _15782_ (.A(_11987_),
    .X(_11990_));
 sky130_fd_sc_hd__a22o_2 _15783_ (.A1(\mem_rdata_q[25] ),
    .A2(_11990_),
    .B1(mem_rdata[25]),
    .B2(_11989_),
    .X(_02956_));
 sky130_fd_sc_hd__a22o_2 _15784_ (.A1(\mem_rdata_q[24] ),
    .A2(_11990_),
    .B1(mem_rdata[24]),
    .B2(_11989_),
    .X(_02955_));
 sky130_fd_sc_hd__a22o_2 _15785_ (.A1(\mem_rdata_q[23] ),
    .A2(_11990_),
    .B1(mem_rdata[23]),
    .B2(_11989_),
    .X(_02954_));
 sky130_fd_sc_hd__a22o_2 _15786_ (.A1(\mem_rdata_q[22] ),
    .A2(_11990_),
    .B1(mem_rdata[22]),
    .B2(_11989_),
    .X(_02953_));
 sky130_fd_sc_hd__buf_1 _15787_ (.A(_10447_),
    .X(_11991_));
 sky130_fd_sc_hd__a22o_2 _15788_ (.A1(\mem_rdata_q[21] ),
    .A2(_11990_),
    .B1(mem_rdata[21]),
    .B2(_11991_),
    .X(_02952_));
 sky130_fd_sc_hd__a22o_2 _15789_ (.A1(\mem_rdata_q[20] ),
    .A2(_11990_),
    .B1(mem_rdata[20]),
    .B2(_11991_),
    .X(_02951_));
 sky130_fd_sc_hd__buf_1 _15790_ (.A(_11987_),
    .X(_11992_));
 sky130_fd_sc_hd__a22o_2 _15791_ (.A1(\mem_rdata_q[19] ),
    .A2(_11992_),
    .B1(mem_rdata[19]),
    .B2(_11991_),
    .X(_02950_));
 sky130_fd_sc_hd__a22o_2 _15792_ (.A1(\mem_rdata_q[18] ),
    .A2(_11992_),
    .B1(mem_rdata[18]),
    .B2(_11991_),
    .X(_02949_));
 sky130_fd_sc_hd__a22o_2 _15793_ (.A1(\mem_rdata_q[17] ),
    .A2(_11992_),
    .B1(mem_rdata[17]),
    .B2(_11991_),
    .X(_02948_));
 sky130_fd_sc_hd__a22o_2 _15794_ (.A1(\mem_rdata_q[16] ),
    .A2(_11992_),
    .B1(mem_rdata[16]),
    .B2(_11991_),
    .X(_02947_));
 sky130_fd_sc_hd__buf_1 _15795_ (.A(_10447_),
    .X(_11993_));
 sky130_fd_sc_hd__a22o_2 _15796_ (.A1(\mem_rdata_q[15] ),
    .A2(_11992_),
    .B1(mem_rdata[15]),
    .B2(_11993_),
    .X(_02946_));
 sky130_fd_sc_hd__a22o_2 _15797_ (.A1(_10727_),
    .A2(_11992_),
    .B1(mem_rdata[14]),
    .B2(_11993_),
    .X(_02945_));
 sky130_fd_sc_hd__buf_1 _15798_ (.A(_11987_),
    .X(_11994_));
 sky130_fd_sc_hd__a22o_2 _15799_ (.A1(_10738_),
    .A2(_11994_),
    .B1(mem_rdata[13]),
    .B2(_11993_),
    .X(_02944_));
 sky130_fd_sc_hd__a22o_2 _15800_ (.A1(_10725_),
    .A2(_11994_),
    .B1(mem_rdata[12]),
    .B2(_11993_),
    .X(_02943_));
 sky130_fd_sc_hd__a22o_2 _15801_ (.A1(\mem_rdata_q[11] ),
    .A2(_11994_),
    .B1(mem_rdata[11]),
    .B2(_11993_),
    .X(_02942_));
 sky130_fd_sc_hd__a22o_2 _15802_ (.A1(\mem_rdata_q[10] ),
    .A2(_11994_),
    .B1(mem_rdata[10]),
    .B2(_11993_),
    .X(_02941_));
 sky130_fd_sc_hd__buf_1 _15803_ (.A(_10447_),
    .X(_11995_));
 sky130_fd_sc_hd__a22o_2 _15804_ (.A1(\mem_rdata_q[9] ),
    .A2(_11994_),
    .B1(mem_rdata[9]),
    .B2(_11995_),
    .X(_02940_));
 sky130_fd_sc_hd__a22o_2 _15805_ (.A1(\mem_rdata_q[8] ),
    .A2(_11994_),
    .B1(mem_rdata[8]),
    .B2(_11995_),
    .X(_02939_));
 sky130_fd_sc_hd__buf_1 _15806_ (.A(_10445_),
    .X(_11996_));
 sky130_fd_sc_hd__a22o_2 _15807_ (.A1(\mem_rdata_q[7] ),
    .A2(_11996_),
    .B1(mem_rdata[7]),
    .B2(_11995_),
    .X(_02938_));
 sky130_fd_sc_hd__a22o_2 _15808_ (.A1(\mem_rdata_q[6] ),
    .A2(_11996_),
    .B1(mem_rdata[6]),
    .B2(_11995_),
    .X(_02937_));
 sky130_fd_sc_hd__a22o_2 _15809_ (.A1(\mem_rdata_q[5] ),
    .A2(_11996_),
    .B1(mem_rdata[5]),
    .B2(_11995_),
    .X(_02936_));
 sky130_fd_sc_hd__a22o_2 _15810_ (.A1(\mem_rdata_q[4] ),
    .A2(_11996_),
    .B1(mem_rdata[4]),
    .B2(_11995_),
    .X(_02935_));
 sky130_fd_sc_hd__a22o_2 _15811_ (.A1(\mem_rdata_q[3] ),
    .A2(_11996_),
    .B1(mem_rdata[3]),
    .B2(_11986_),
    .X(_02934_));
 sky130_fd_sc_hd__a22o_2 _15812_ (.A1(\mem_rdata_q[2] ),
    .A2(_11996_),
    .B1(mem_rdata[2]),
    .B2(_11986_),
    .X(_02933_));
 sky130_fd_sc_hd__a22o_2 _15813_ (.A1(\mem_rdata_q[1] ),
    .A2(_11987_),
    .B1(mem_rdata[1]),
    .B2(_11986_),
    .X(_02932_));
 sky130_fd_sc_hd__a22o_2 _15814_ (.A1(\mem_rdata_q[0] ),
    .A2(_11987_),
    .B1(mem_rdata[0]),
    .B2(_11986_),
    .X(_02931_));
 sky130_fd_sc_hd__or4_2 _15815_ (.A(_11380_),
    .B(_11310_),
    .C(_11252_),
    .D(_11262_),
    .X(_11997_));
 sky130_fd_sc_hd__buf_1 _15816_ (.A(_11997_),
    .X(_11998_));
 sky130_fd_sc_hd__buf_1 _15817_ (.A(_11998_),
    .X(_11999_));
 sky130_vsdinv _15818_ (.A(_11997_),
    .Y(_12000_));
 sky130_fd_sc_hd__buf_1 _15819_ (.A(_12000_),
    .X(_12001_));
 sky130_fd_sc_hd__buf_1 _15820_ (.A(_12001_),
    .X(_12002_));
 sky130_fd_sc_hd__a22o_2 _15821_ (.A1(\cpuregs[18][31] ),
    .A2(_11999_),
    .B1(_11653_),
    .B2(_12002_),
    .X(_02930_));
 sky130_fd_sc_hd__a22o_2 _15822_ (.A1(\cpuregs[18][30] ),
    .A2(_11999_),
    .B1(_11657_),
    .B2(_12002_),
    .X(_02929_));
 sky130_fd_sc_hd__a22o_2 _15823_ (.A1(\cpuregs[18][29] ),
    .A2(_11999_),
    .B1(_11658_),
    .B2(_12002_),
    .X(_02928_));
 sky130_fd_sc_hd__a22o_2 _15824_ (.A1(\cpuregs[18][28] ),
    .A2(_11999_),
    .B1(_11659_),
    .B2(_12002_),
    .X(_02927_));
 sky130_fd_sc_hd__a22o_2 _15825_ (.A1(\cpuregs[18][27] ),
    .A2(_11999_),
    .B1(_11660_),
    .B2(_12002_),
    .X(_02926_));
 sky130_fd_sc_hd__a22o_2 _15826_ (.A1(\cpuregs[18][26] ),
    .A2(_11999_),
    .B1(_11661_),
    .B2(_12002_),
    .X(_02925_));
 sky130_fd_sc_hd__buf_1 _15827_ (.A(_11998_),
    .X(_12003_));
 sky130_fd_sc_hd__buf_1 _15828_ (.A(_12001_),
    .X(_12004_));
 sky130_fd_sc_hd__a22o_2 _15829_ (.A1(\cpuregs[18][25] ),
    .A2(_12003_),
    .B1(_11663_),
    .B2(_12004_),
    .X(_02924_));
 sky130_fd_sc_hd__a22o_2 _15830_ (.A1(\cpuregs[18][24] ),
    .A2(_12003_),
    .B1(_11665_),
    .B2(_12004_),
    .X(_02923_));
 sky130_fd_sc_hd__a22o_2 _15831_ (.A1(\cpuregs[18][23] ),
    .A2(_12003_),
    .B1(_11666_),
    .B2(_12004_),
    .X(_02922_));
 sky130_fd_sc_hd__a22o_2 _15832_ (.A1(\cpuregs[18][22] ),
    .A2(_12003_),
    .B1(_11667_),
    .B2(_12004_),
    .X(_02921_));
 sky130_fd_sc_hd__a22o_2 _15833_ (.A1(\cpuregs[18][21] ),
    .A2(_12003_),
    .B1(_11668_),
    .B2(_12004_),
    .X(_02920_));
 sky130_fd_sc_hd__a22o_2 _15834_ (.A1(\cpuregs[18][20] ),
    .A2(_12003_),
    .B1(_11669_),
    .B2(_12004_),
    .X(_02919_));
 sky130_fd_sc_hd__buf_1 _15835_ (.A(_11998_),
    .X(_12005_));
 sky130_fd_sc_hd__buf_1 _15836_ (.A(_12001_),
    .X(_12006_));
 sky130_fd_sc_hd__a22o_2 _15837_ (.A1(\cpuregs[18][19] ),
    .A2(_12005_),
    .B1(_11671_),
    .B2(_12006_),
    .X(_02918_));
 sky130_fd_sc_hd__a22o_2 _15838_ (.A1(\cpuregs[18][18] ),
    .A2(_12005_),
    .B1(_11673_),
    .B2(_12006_),
    .X(_02917_));
 sky130_fd_sc_hd__a22o_2 _15839_ (.A1(\cpuregs[18][17] ),
    .A2(_12005_),
    .B1(_11674_),
    .B2(_12006_),
    .X(_02916_));
 sky130_fd_sc_hd__a22o_2 _15840_ (.A1(\cpuregs[18][16] ),
    .A2(_12005_),
    .B1(_11675_),
    .B2(_12006_),
    .X(_02915_));
 sky130_fd_sc_hd__a22o_2 _15841_ (.A1(\cpuregs[18][15] ),
    .A2(_12005_),
    .B1(_11676_),
    .B2(_12006_),
    .X(_02914_));
 sky130_fd_sc_hd__a22o_2 _15842_ (.A1(\cpuregs[18][14] ),
    .A2(_12005_),
    .B1(_11677_),
    .B2(_12006_),
    .X(_02913_));
 sky130_fd_sc_hd__buf_1 _15843_ (.A(_11998_),
    .X(_12007_));
 sky130_fd_sc_hd__buf_1 _15844_ (.A(_12001_),
    .X(_12008_));
 sky130_fd_sc_hd__a22o_2 _15845_ (.A1(\cpuregs[18][13] ),
    .A2(_12007_),
    .B1(_11679_),
    .B2(_12008_),
    .X(_02912_));
 sky130_fd_sc_hd__a22o_2 _15846_ (.A1(\cpuregs[18][12] ),
    .A2(_12007_),
    .B1(_11681_),
    .B2(_12008_),
    .X(_02911_));
 sky130_fd_sc_hd__a22o_2 _15847_ (.A1(\cpuregs[18][11] ),
    .A2(_12007_),
    .B1(_11682_),
    .B2(_12008_),
    .X(_02910_));
 sky130_fd_sc_hd__a22o_2 _15848_ (.A1(\cpuregs[18][10] ),
    .A2(_12007_),
    .B1(_11683_),
    .B2(_12008_),
    .X(_02909_));
 sky130_fd_sc_hd__a22o_2 _15849_ (.A1(\cpuregs[18][9] ),
    .A2(_12007_),
    .B1(_11684_),
    .B2(_12008_),
    .X(_02908_));
 sky130_fd_sc_hd__a22o_2 _15850_ (.A1(\cpuregs[18][8] ),
    .A2(_12007_),
    .B1(_11685_),
    .B2(_12008_),
    .X(_02907_));
 sky130_fd_sc_hd__buf_1 _15851_ (.A(_11997_),
    .X(_12009_));
 sky130_fd_sc_hd__buf_1 _15852_ (.A(_12000_),
    .X(_12010_));
 sky130_fd_sc_hd__a22o_2 _15853_ (.A1(\cpuregs[18][7] ),
    .A2(_12009_),
    .B1(_11687_),
    .B2(_12010_),
    .X(_02906_));
 sky130_fd_sc_hd__a22o_2 _15854_ (.A1(\cpuregs[18][6] ),
    .A2(_12009_),
    .B1(_11689_),
    .B2(_12010_),
    .X(_02905_));
 sky130_fd_sc_hd__a22o_2 _15855_ (.A1(\cpuregs[18][5] ),
    .A2(_12009_),
    .B1(_11690_),
    .B2(_12010_),
    .X(_02904_));
 sky130_fd_sc_hd__a22o_2 _15856_ (.A1(\cpuregs[18][4] ),
    .A2(_12009_),
    .B1(_11691_),
    .B2(_12010_),
    .X(_02903_));
 sky130_fd_sc_hd__a22o_2 _15857_ (.A1(\cpuregs[18][3] ),
    .A2(_12009_),
    .B1(_11692_),
    .B2(_12010_),
    .X(_02902_));
 sky130_fd_sc_hd__a22o_2 _15858_ (.A1(\cpuregs[18][2] ),
    .A2(_12009_),
    .B1(_11693_),
    .B2(_12010_),
    .X(_02901_));
 sky130_fd_sc_hd__a22o_2 _15859_ (.A1(\cpuregs[18][1] ),
    .A2(_11998_),
    .B1(_11694_),
    .B2(_12001_),
    .X(_02900_));
 sky130_fd_sc_hd__a22o_2 _15860_ (.A1(\cpuregs[18][0] ),
    .A2(_11998_),
    .B1(_11695_),
    .B2(_12001_),
    .X(_02899_));
 sky130_fd_sc_hd__or2_2 _15861_ (.A(_11262_),
    .B(_11311_),
    .X(_12011_));
 sky130_fd_sc_hd__buf_1 _15862_ (.A(_12011_),
    .X(_12012_));
 sky130_fd_sc_hd__buf_1 _15863_ (.A(_12012_),
    .X(_12013_));
 sky130_vsdinv _15864_ (.A(_12011_),
    .Y(_12014_));
 sky130_fd_sc_hd__buf_1 _15865_ (.A(_12014_),
    .X(_12015_));
 sky130_fd_sc_hd__buf_1 _15866_ (.A(_12015_),
    .X(_12016_));
 sky130_fd_sc_hd__a22o_2 _15867_ (.A1(\cpuregs[10][31] ),
    .A2(_12013_),
    .B1(_11653_),
    .B2(_12016_),
    .X(_02898_));
 sky130_fd_sc_hd__a22o_2 _15868_ (.A1(\cpuregs[10][30] ),
    .A2(_12013_),
    .B1(_11657_),
    .B2(_12016_),
    .X(_02897_));
 sky130_fd_sc_hd__a22o_2 _15869_ (.A1(\cpuregs[10][29] ),
    .A2(_12013_),
    .B1(_11658_),
    .B2(_12016_),
    .X(_02896_));
 sky130_fd_sc_hd__a22o_2 _15870_ (.A1(\cpuregs[10][28] ),
    .A2(_12013_),
    .B1(_11659_),
    .B2(_12016_),
    .X(_02895_));
 sky130_fd_sc_hd__a22o_2 _15871_ (.A1(\cpuregs[10][27] ),
    .A2(_12013_),
    .B1(_11660_),
    .B2(_12016_),
    .X(_02894_));
 sky130_fd_sc_hd__a22o_2 _15872_ (.A1(\cpuregs[10][26] ),
    .A2(_12013_),
    .B1(_11661_),
    .B2(_12016_),
    .X(_02893_));
 sky130_fd_sc_hd__buf_1 _15873_ (.A(_12012_),
    .X(_12017_));
 sky130_fd_sc_hd__buf_1 _15874_ (.A(_12015_),
    .X(_12018_));
 sky130_fd_sc_hd__a22o_2 _15875_ (.A1(\cpuregs[10][25] ),
    .A2(_12017_),
    .B1(_11663_),
    .B2(_12018_),
    .X(_02892_));
 sky130_fd_sc_hd__a22o_2 _15876_ (.A1(\cpuregs[10][24] ),
    .A2(_12017_),
    .B1(_11665_),
    .B2(_12018_),
    .X(_02891_));
 sky130_fd_sc_hd__a22o_2 _15877_ (.A1(\cpuregs[10][23] ),
    .A2(_12017_),
    .B1(_11666_),
    .B2(_12018_),
    .X(_02890_));
 sky130_fd_sc_hd__a22o_2 _15878_ (.A1(\cpuregs[10][22] ),
    .A2(_12017_),
    .B1(_11667_),
    .B2(_12018_),
    .X(_02889_));
 sky130_fd_sc_hd__a22o_2 _15879_ (.A1(\cpuregs[10][21] ),
    .A2(_12017_),
    .B1(_11668_),
    .B2(_12018_),
    .X(_02888_));
 sky130_fd_sc_hd__a22o_2 _15880_ (.A1(\cpuregs[10][20] ),
    .A2(_12017_),
    .B1(_11669_),
    .B2(_12018_),
    .X(_02887_));
 sky130_fd_sc_hd__buf_1 _15881_ (.A(_12012_),
    .X(_12019_));
 sky130_fd_sc_hd__buf_1 _15882_ (.A(_12015_),
    .X(_12020_));
 sky130_fd_sc_hd__a22o_2 _15883_ (.A1(\cpuregs[10][19] ),
    .A2(_12019_),
    .B1(_11671_),
    .B2(_12020_),
    .X(_02886_));
 sky130_fd_sc_hd__a22o_2 _15884_ (.A1(\cpuregs[10][18] ),
    .A2(_12019_),
    .B1(_11673_),
    .B2(_12020_),
    .X(_02885_));
 sky130_fd_sc_hd__a22o_2 _15885_ (.A1(\cpuregs[10][17] ),
    .A2(_12019_),
    .B1(_11674_),
    .B2(_12020_),
    .X(_02884_));
 sky130_fd_sc_hd__a22o_2 _15886_ (.A1(\cpuregs[10][16] ),
    .A2(_12019_),
    .B1(_11675_),
    .B2(_12020_),
    .X(_02883_));
 sky130_fd_sc_hd__a22o_2 _15887_ (.A1(\cpuregs[10][15] ),
    .A2(_12019_),
    .B1(_11676_),
    .B2(_12020_),
    .X(_02882_));
 sky130_fd_sc_hd__a22o_2 _15888_ (.A1(\cpuregs[10][14] ),
    .A2(_12019_),
    .B1(_11677_),
    .B2(_12020_),
    .X(_02881_));
 sky130_fd_sc_hd__buf_1 _15889_ (.A(_12012_),
    .X(_12021_));
 sky130_fd_sc_hd__buf_1 _15890_ (.A(_12015_),
    .X(_12022_));
 sky130_fd_sc_hd__a22o_2 _15891_ (.A1(\cpuregs[10][13] ),
    .A2(_12021_),
    .B1(_11679_),
    .B2(_12022_),
    .X(_02880_));
 sky130_fd_sc_hd__a22o_2 _15892_ (.A1(\cpuregs[10][12] ),
    .A2(_12021_),
    .B1(_11681_),
    .B2(_12022_),
    .X(_02879_));
 sky130_fd_sc_hd__a22o_2 _15893_ (.A1(\cpuregs[10][11] ),
    .A2(_12021_),
    .B1(_11682_),
    .B2(_12022_),
    .X(_02878_));
 sky130_fd_sc_hd__a22o_2 _15894_ (.A1(\cpuregs[10][10] ),
    .A2(_12021_),
    .B1(_11683_),
    .B2(_12022_),
    .X(_02877_));
 sky130_fd_sc_hd__a22o_2 _15895_ (.A1(\cpuregs[10][9] ),
    .A2(_12021_),
    .B1(_11684_),
    .B2(_12022_),
    .X(_02876_));
 sky130_fd_sc_hd__a22o_2 _15896_ (.A1(\cpuregs[10][8] ),
    .A2(_12021_),
    .B1(_11685_),
    .B2(_12022_),
    .X(_02875_));
 sky130_fd_sc_hd__buf_1 _15897_ (.A(_12011_),
    .X(_12023_));
 sky130_fd_sc_hd__buf_1 _15898_ (.A(_12014_),
    .X(_12024_));
 sky130_fd_sc_hd__a22o_2 _15899_ (.A1(\cpuregs[10][7] ),
    .A2(_12023_),
    .B1(_11687_),
    .B2(_12024_),
    .X(_02874_));
 sky130_fd_sc_hd__a22o_2 _15900_ (.A1(\cpuregs[10][6] ),
    .A2(_12023_),
    .B1(_11689_),
    .B2(_12024_),
    .X(_02873_));
 sky130_fd_sc_hd__a22o_2 _15901_ (.A1(\cpuregs[10][5] ),
    .A2(_12023_),
    .B1(_11690_),
    .B2(_12024_),
    .X(_02872_));
 sky130_fd_sc_hd__a22o_2 _15902_ (.A1(\cpuregs[10][4] ),
    .A2(_12023_),
    .B1(_11691_),
    .B2(_12024_),
    .X(_02871_));
 sky130_fd_sc_hd__a22o_2 _15903_ (.A1(\cpuregs[10][3] ),
    .A2(_12023_),
    .B1(_11692_),
    .B2(_12024_),
    .X(_02870_));
 sky130_fd_sc_hd__a22o_2 _15904_ (.A1(\cpuregs[10][2] ),
    .A2(_12023_),
    .B1(_11693_),
    .B2(_12024_),
    .X(_02869_));
 sky130_fd_sc_hd__a22o_2 _15905_ (.A1(\cpuregs[10][1] ),
    .A2(_12012_),
    .B1(_11694_),
    .B2(_12015_),
    .X(_02868_));
 sky130_fd_sc_hd__a22o_2 _15906_ (.A1(\cpuregs[10][0] ),
    .A2(_12012_),
    .B1(_11695_),
    .B2(_12015_),
    .X(_02867_));
 sky130_fd_sc_hd__buf_1 _15907_ (.A(\cpuregs[0][31] ),
    .X(_02866_));
 sky130_fd_sc_hd__buf_1 _15908_ (.A(\cpuregs[0][30] ),
    .X(_02865_));
 sky130_fd_sc_hd__buf_1 _15909_ (.A(\cpuregs[0][29] ),
    .X(_02864_));
 sky130_fd_sc_hd__buf_1 _15910_ (.A(\cpuregs[0][28] ),
    .X(_02863_));
 sky130_fd_sc_hd__buf_1 _15911_ (.A(\cpuregs[0][27] ),
    .X(_02862_));
 sky130_fd_sc_hd__buf_1 _15912_ (.A(\cpuregs[0][26] ),
    .X(_02861_));
 sky130_fd_sc_hd__buf_1 _15913_ (.A(\cpuregs[0][25] ),
    .X(_02860_));
 sky130_fd_sc_hd__buf_1 _15914_ (.A(\cpuregs[0][24] ),
    .X(_02859_));
 sky130_fd_sc_hd__buf_1 _15915_ (.A(\cpuregs[0][23] ),
    .X(_02858_));
 sky130_fd_sc_hd__buf_1 _15916_ (.A(\cpuregs[0][22] ),
    .X(_02857_));
 sky130_fd_sc_hd__buf_1 _15917_ (.A(\cpuregs[0][21] ),
    .X(_02856_));
 sky130_fd_sc_hd__buf_1 _15918_ (.A(\cpuregs[0][20] ),
    .X(_02855_));
 sky130_fd_sc_hd__buf_1 _15919_ (.A(\cpuregs[0][19] ),
    .X(_02854_));
 sky130_fd_sc_hd__buf_1 _15920_ (.A(\cpuregs[0][18] ),
    .X(_02853_));
 sky130_fd_sc_hd__buf_1 _15921_ (.A(\cpuregs[0][17] ),
    .X(_02852_));
 sky130_fd_sc_hd__buf_1 _15922_ (.A(\cpuregs[0][16] ),
    .X(_02851_));
 sky130_fd_sc_hd__buf_1 _15923_ (.A(\cpuregs[0][15] ),
    .X(_02850_));
 sky130_fd_sc_hd__buf_1 _15924_ (.A(\cpuregs[0][14] ),
    .X(_02849_));
 sky130_fd_sc_hd__buf_1 _15925_ (.A(\cpuregs[0][13] ),
    .X(_02848_));
 sky130_fd_sc_hd__buf_1 _15926_ (.A(\cpuregs[0][12] ),
    .X(_02847_));
 sky130_fd_sc_hd__buf_1 _15927_ (.A(\cpuregs[0][11] ),
    .X(_02846_));
 sky130_fd_sc_hd__buf_1 _15928_ (.A(\cpuregs[0][10] ),
    .X(_02845_));
 sky130_fd_sc_hd__buf_1 _15929_ (.A(\cpuregs[0][9] ),
    .X(_02844_));
 sky130_fd_sc_hd__buf_1 _15930_ (.A(\cpuregs[0][8] ),
    .X(_02843_));
 sky130_fd_sc_hd__buf_1 _15931_ (.A(\cpuregs[0][7] ),
    .X(_02842_));
 sky130_fd_sc_hd__buf_1 _15932_ (.A(\cpuregs[0][6] ),
    .X(_02841_));
 sky130_fd_sc_hd__buf_1 _15933_ (.A(\cpuregs[0][5] ),
    .X(_02840_));
 sky130_fd_sc_hd__buf_1 _15934_ (.A(\cpuregs[0][4] ),
    .X(_02839_));
 sky130_fd_sc_hd__buf_1 _15935_ (.A(\cpuregs[0][3] ),
    .X(_02838_));
 sky130_fd_sc_hd__buf_1 _15936_ (.A(\cpuregs[0][2] ),
    .X(_02837_));
 sky130_fd_sc_hd__buf_1 _15937_ (.A(\cpuregs[0][1] ),
    .X(_02836_));
 sky130_fd_sc_hd__buf_1 _15938_ (.A(\cpuregs[0][0] ),
    .X(_02835_));
 sky130_fd_sc_hd__or2_2 _15939_ (.A(_11262_),
    .B(_11428_),
    .X(_12025_));
 sky130_fd_sc_hd__buf_1 _15940_ (.A(_12025_),
    .X(_12026_));
 sky130_fd_sc_hd__buf_1 _15941_ (.A(_12026_),
    .X(_12027_));
 sky130_vsdinv _15942_ (.A(_12025_),
    .Y(_12028_));
 sky130_fd_sc_hd__buf_1 _15943_ (.A(_12028_),
    .X(_12029_));
 sky130_fd_sc_hd__buf_1 _15944_ (.A(_12029_),
    .X(_12030_));
 sky130_fd_sc_hd__a22o_2 _15945_ (.A1(\cpuregs[14][31] ),
    .A2(_12027_),
    .B1(_11653_),
    .B2(_12030_),
    .X(_02834_));
 sky130_fd_sc_hd__a22o_2 _15946_ (.A1(\cpuregs[14][30] ),
    .A2(_12027_),
    .B1(_11657_),
    .B2(_12030_),
    .X(_02833_));
 sky130_fd_sc_hd__a22o_2 _15947_ (.A1(\cpuregs[14][29] ),
    .A2(_12027_),
    .B1(_11658_),
    .B2(_12030_),
    .X(_02832_));
 sky130_fd_sc_hd__a22o_2 _15948_ (.A1(\cpuregs[14][28] ),
    .A2(_12027_),
    .B1(_11659_),
    .B2(_12030_),
    .X(_02831_));
 sky130_fd_sc_hd__a22o_2 _15949_ (.A1(\cpuregs[14][27] ),
    .A2(_12027_),
    .B1(_11660_),
    .B2(_12030_),
    .X(_02830_));
 sky130_fd_sc_hd__a22o_2 _15950_ (.A1(\cpuregs[14][26] ),
    .A2(_12027_),
    .B1(_11661_),
    .B2(_12030_),
    .X(_02829_));
 sky130_fd_sc_hd__buf_1 _15951_ (.A(_12026_),
    .X(_12031_));
 sky130_fd_sc_hd__buf_1 _15952_ (.A(_12029_),
    .X(_12032_));
 sky130_fd_sc_hd__a22o_2 _15953_ (.A1(\cpuregs[14][25] ),
    .A2(_12031_),
    .B1(_11663_),
    .B2(_12032_),
    .X(_02828_));
 sky130_fd_sc_hd__a22o_2 _15954_ (.A1(\cpuregs[14][24] ),
    .A2(_12031_),
    .B1(_11665_),
    .B2(_12032_),
    .X(_02827_));
 sky130_fd_sc_hd__a22o_2 _15955_ (.A1(\cpuregs[14][23] ),
    .A2(_12031_),
    .B1(_11666_),
    .B2(_12032_),
    .X(_02826_));
 sky130_fd_sc_hd__a22o_2 _15956_ (.A1(\cpuregs[14][22] ),
    .A2(_12031_),
    .B1(_11667_),
    .B2(_12032_),
    .X(_02825_));
 sky130_fd_sc_hd__a22o_2 _15957_ (.A1(\cpuregs[14][21] ),
    .A2(_12031_),
    .B1(_11668_),
    .B2(_12032_),
    .X(_02824_));
 sky130_fd_sc_hd__a22o_2 _15958_ (.A1(\cpuregs[14][20] ),
    .A2(_12031_),
    .B1(_11669_),
    .B2(_12032_),
    .X(_02823_));
 sky130_fd_sc_hd__buf_1 _15959_ (.A(_12026_),
    .X(_12033_));
 sky130_fd_sc_hd__buf_1 _15960_ (.A(_12029_),
    .X(_12034_));
 sky130_fd_sc_hd__a22o_2 _15961_ (.A1(\cpuregs[14][19] ),
    .A2(_12033_),
    .B1(_11671_),
    .B2(_12034_),
    .X(_02822_));
 sky130_fd_sc_hd__a22o_2 _15962_ (.A1(\cpuregs[14][18] ),
    .A2(_12033_),
    .B1(_11673_),
    .B2(_12034_),
    .X(_02821_));
 sky130_fd_sc_hd__a22o_2 _15963_ (.A1(\cpuregs[14][17] ),
    .A2(_12033_),
    .B1(_11674_),
    .B2(_12034_),
    .X(_02820_));
 sky130_fd_sc_hd__a22o_2 _15964_ (.A1(\cpuregs[14][16] ),
    .A2(_12033_),
    .B1(_11675_),
    .B2(_12034_),
    .X(_02819_));
 sky130_fd_sc_hd__a22o_2 _15965_ (.A1(\cpuregs[14][15] ),
    .A2(_12033_),
    .B1(_11676_),
    .B2(_12034_),
    .X(_02818_));
 sky130_fd_sc_hd__a22o_2 _15966_ (.A1(\cpuregs[14][14] ),
    .A2(_12033_),
    .B1(_11677_),
    .B2(_12034_),
    .X(_02817_));
 sky130_fd_sc_hd__buf_1 _15967_ (.A(_12026_),
    .X(_12035_));
 sky130_fd_sc_hd__buf_1 _15968_ (.A(_12029_),
    .X(_12036_));
 sky130_fd_sc_hd__a22o_2 _15969_ (.A1(\cpuregs[14][13] ),
    .A2(_12035_),
    .B1(_11679_),
    .B2(_12036_),
    .X(_02816_));
 sky130_fd_sc_hd__a22o_2 _15970_ (.A1(\cpuregs[14][12] ),
    .A2(_12035_),
    .B1(_11681_),
    .B2(_12036_),
    .X(_02815_));
 sky130_fd_sc_hd__a22o_2 _15971_ (.A1(\cpuregs[14][11] ),
    .A2(_12035_),
    .B1(_11682_),
    .B2(_12036_),
    .X(_02814_));
 sky130_fd_sc_hd__a22o_2 _15972_ (.A1(\cpuregs[14][10] ),
    .A2(_12035_),
    .B1(_11683_),
    .B2(_12036_),
    .X(_02813_));
 sky130_fd_sc_hd__a22o_2 _15973_ (.A1(\cpuregs[14][9] ),
    .A2(_12035_),
    .B1(_11684_),
    .B2(_12036_),
    .X(_02812_));
 sky130_fd_sc_hd__a22o_2 _15974_ (.A1(\cpuregs[14][8] ),
    .A2(_12035_),
    .B1(_11685_),
    .B2(_12036_),
    .X(_02811_));
 sky130_fd_sc_hd__buf_1 _15975_ (.A(_12025_),
    .X(_12037_));
 sky130_fd_sc_hd__buf_1 _15976_ (.A(_12028_),
    .X(_12038_));
 sky130_fd_sc_hd__a22o_2 _15977_ (.A1(\cpuregs[14][7] ),
    .A2(_12037_),
    .B1(_11687_),
    .B2(_12038_),
    .X(_02810_));
 sky130_fd_sc_hd__a22o_2 _15978_ (.A1(\cpuregs[14][6] ),
    .A2(_12037_),
    .B1(_11689_),
    .B2(_12038_),
    .X(_02809_));
 sky130_fd_sc_hd__a22o_2 _15979_ (.A1(\cpuregs[14][5] ),
    .A2(_12037_),
    .B1(_11690_),
    .B2(_12038_),
    .X(_02808_));
 sky130_fd_sc_hd__a22o_2 _15980_ (.A1(\cpuregs[14][4] ),
    .A2(_12037_),
    .B1(_11691_),
    .B2(_12038_),
    .X(_02807_));
 sky130_fd_sc_hd__a22o_2 _15981_ (.A1(\cpuregs[14][3] ),
    .A2(_12037_),
    .B1(_11692_),
    .B2(_12038_),
    .X(_02806_));
 sky130_fd_sc_hd__a22o_2 _15982_ (.A1(\cpuregs[14][2] ),
    .A2(_12037_),
    .B1(_11693_),
    .B2(_12038_),
    .X(_02805_));
 sky130_fd_sc_hd__a22o_2 _15983_ (.A1(\cpuregs[14][1] ),
    .A2(_12026_),
    .B1(_11694_),
    .B2(_12029_),
    .X(_02804_));
 sky130_fd_sc_hd__a22o_2 _15984_ (.A1(\cpuregs[14][0] ),
    .A2(_12026_),
    .B1(_11695_),
    .B2(_12029_),
    .X(_02803_));
 sky130_fd_sc_hd__or2_2 _15985_ (.A(_11311_),
    .B(_11365_),
    .X(_12039_));
 sky130_fd_sc_hd__buf_1 _15986_ (.A(_12039_),
    .X(_12040_));
 sky130_fd_sc_hd__buf_1 _15987_ (.A(_12040_),
    .X(_12041_));
 sky130_vsdinv _15988_ (.A(_12039_),
    .Y(_12042_));
 sky130_fd_sc_hd__buf_1 _15989_ (.A(_12042_),
    .X(_12043_));
 sky130_fd_sc_hd__buf_1 _15990_ (.A(_12043_),
    .X(_12044_));
 sky130_fd_sc_hd__a22o_2 _15991_ (.A1(\cpuregs[8][31] ),
    .A2(_12041_),
    .B1(\cpuregs_wrdata[31] ),
    .B2(_12044_),
    .X(_02802_));
 sky130_fd_sc_hd__a22o_2 _15992_ (.A1(\cpuregs[8][30] ),
    .A2(_12041_),
    .B1(\cpuregs_wrdata[30] ),
    .B2(_12044_),
    .X(_02801_));
 sky130_fd_sc_hd__a22o_2 _15993_ (.A1(\cpuregs[8][29] ),
    .A2(_12041_),
    .B1(\cpuregs_wrdata[29] ),
    .B2(_12044_),
    .X(_02800_));
 sky130_fd_sc_hd__a22o_2 _15994_ (.A1(\cpuregs[8][28] ),
    .A2(_12041_),
    .B1(\cpuregs_wrdata[28] ),
    .B2(_12044_),
    .X(_02799_));
 sky130_fd_sc_hd__a22o_2 _15995_ (.A1(\cpuregs[8][27] ),
    .A2(_12041_),
    .B1(\cpuregs_wrdata[27] ),
    .B2(_12044_),
    .X(_02798_));
 sky130_fd_sc_hd__a22o_2 _15996_ (.A1(\cpuregs[8][26] ),
    .A2(_12041_),
    .B1(\cpuregs_wrdata[26] ),
    .B2(_12044_),
    .X(_02797_));
 sky130_fd_sc_hd__buf_1 _15997_ (.A(_12040_),
    .X(_12045_));
 sky130_fd_sc_hd__buf_1 _15998_ (.A(_12043_),
    .X(_12046_));
 sky130_fd_sc_hd__a22o_2 _15999_ (.A1(\cpuregs[8][25] ),
    .A2(_12045_),
    .B1(\cpuregs_wrdata[25] ),
    .B2(_12046_),
    .X(_02796_));
 sky130_fd_sc_hd__a22o_2 _16000_ (.A1(\cpuregs[8][24] ),
    .A2(_12045_),
    .B1(\cpuregs_wrdata[24] ),
    .B2(_12046_),
    .X(_02795_));
 sky130_fd_sc_hd__a22o_2 _16001_ (.A1(\cpuregs[8][23] ),
    .A2(_12045_),
    .B1(\cpuregs_wrdata[23] ),
    .B2(_12046_),
    .X(_02794_));
 sky130_fd_sc_hd__a22o_2 _16002_ (.A1(\cpuregs[8][22] ),
    .A2(_12045_),
    .B1(\cpuregs_wrdata[22] ),
    .B2(_12046_),
    .X(_02793_));
 sky130_fd_sc_hd__a22o_2 _16003_ (.A1(\cpuregs[8][21] ),
    .A2(_12045_),
    .B1(\cpuregs_wrdata[21] ),
    .B2(_12046_),
    .X(_02792_));
 sky130_fd_sc_hd__a22o_2 _16004_ (.A1(\cpuregs[8][20] ),
    .A2(_12045_),
    .B1(\cpuregs_wrdata[20] ),
    .B2(_12046_),
    .X(_02791_));
 sky130_fd_sc_hd__buf_1 _16005_ (.A(_12040_),
    .X(_12047_));
 sky130_fd_sc_hd__buf_1 _16006_ (.A(_12043_),
    .X(_12048_));
 sky130_fd_sc_hd__a22o_2 _16007_ (.A1(\cpuregs[8][19] ),
    .A2(_12047_),
    .B1(\cpuregs_wrdata[19] ),
    .B2(_12048_),
    .X(_02790_));
 sky130_fd_sc_hd__a22o_2 _16008_ (.A1(\cpuregs[8][18] ),
    .A2(_12047_),
    .B1(\cpuregs_wrdata[18] ),
    .B2(_12048_),
    .X(_02789_));
 sky130_fd_sc_hd__a22o_2 _16009_ (.A1(\cpuregs[8][17] ),
    .A2(_12047_),
    .B1(\cpuregs_wrdata[17] ),
    .B2(_12048_),
    .X(_02788_));
 sky130_fd_sc_hd__a22o_2 _16010_ (.A1(\cpuregs[8][16] ),
    .A2(_12047_),
    .B1(\cpuregs_wrdata[16] ),
    .B2(_12048_),
    .X(_02787_));
 sky130_fd_sc_hd__a22o_2 _16011_ (.A1(\cpuregs[8][15] ),
    .A2(_12047_),
    .B1(\cpuregs_wrdata[15] ),
    .B2(_12048_),
    .X(_02786_));
 sky130_fd_sc_hd__a22o_2 _16012_ (.A1(\cpuregs[8][14] ),
    .A2(_12047_),
    .B1(\cpuregs_wrdata[14] ),
    .B2(_12048_),
    .X(_02785_));
 sky130_fd_sc_hd__buf_1 _16013_ (.A(_12040_),
    .X(_12049_));
 sky130_fd_sc_hd__buf_1 _16014_ (.A(_12043_),
    .X(_12050_));
 sky130_fd_sc_hd__a22o_2 _16015_ (.A1(\cpuregs[8][13] ),
    .A2(_12049_),
    .B1(\cpuregs_wrdata[13] ),
    .B2(_12050_),
    .X(_02784_));
 sky130_fd_sc_hd__a22o_2 _16016_ (.A1(\cpuregs[8][12] ),
    .A2(_12049_),
    .B1(\cpuregs_wrdata[12] ),
    .B2(_12050_),
    .X(_02783_));
 sky130_fd_sc_hd__a22o_2 _16017_ (.A1(\cpuregs[8][11] ),
    .A2(_12049_),
    .B1(\cpuregs_wrdata[11] ),
    .B2(_12050_),
    .X(_02782_));
 sky130_fd_sc_hd__a22o_2 _16018_ (.A1(\cpuregs[8][10] ),
    .A2(_12049_),
    .B1(\cpuregs_wrdata[10] ),
    .B2(_12050_),
    .X(_02781_));
 sky130_fd_sc_hd__a22o_2 _16019_ (.A1(\cpuregs[8][9] ),
    .A2(_12049_),
    .B1(\cpuregs_wrdata[9] ),
    .B2(_12050_),
    .X(_02780_));
 sky130_fd_sc_hd__a22o_2 _16020_ (.A1(\cpuregs[8][8] ),
    .A2(_12049_),
    .B1(\cpuregs_wrdata[8] ),
    .B2(_12050_),
    .X(_02779_));
 sky130_fd_sc_hd__buf_1 _16021_ (.A(_12039_),
    .X(_12051_));
 sky130_fd_sc_hd__buf_1 _16022_ (.A(_12042_),
    .X(_12052_));
 sky130_fd_sc_hd__a22o_2 _16023_ (.A1(\cpuregs[8][7] ),
    .A2(_12051_),
    .B1(\cpuregs_wrdata[7] ),
    .B2(_12052_),
    .X(_02778_));
 sky130_fd_sc_hd__a22o_2 _16024_ (.A1(\cpuregs[8][6] ),
    .A2(_12051_),
    .B1(\cpuregs_wrdata[6] ),
    .B2(_12052_),
    .X(_02777_));
 sky130_fd_sc_hd__a22o_2 _16025_ (.A1(\cpuregs[8][5] ),
    .A2(_12051_),
    .B1(\cpuregs_wrdata[5] ),
    .B2(_12052_),
    .X(_02776_));
 sky130_fd_sc_hd__a22o_2 _16026_ (.A1(\cpuregs[8][4] ),
    .A2(_12051_),
    .B1(\cpuregs_wrdata[4] ),
    .B2(_12052_),
    .X(_02775_));
 sky130_fd_sc_hd__a22o_2 _16027_ (.A1(\cpuregs[8][3] ),
    .A2(_12051_),
    .B1(\cpuregs_wrdata[3] ),
    .B2(_12052_),
    .X(_02774_));
 sky130_fd_sc_hd__a22o_2 _16028_ (.A1(\cpuregs[8][2] ),
    .A2(_12051_),
    .B1(\cpuregs_wrdata[2] ),
    .B2(_12052_),
    .X(_02773_));
 sky130_fd_sc_hd__a22o_2 _16029_ (.A1(\cpuregs[8][1] ),
    .A2(_12040_),
    .B1(\cpuregs_wrdata[1] ),
    .B2(_12043_),
    .X(_02772_));
 sky130_fd_sc_hd__a22o_2 _16030_ (.A1(\cpuregs[8][0] ),
    .A2(_12040_),
    .B1(\cpuregs_wrdata[0] ),
    .B2(_12043_),
    .X(_02771_));
 sky130_fd_sc_hd__nor2_2 _16031_ (.A(latched_branch),
    .B(_10655_),
    .Y(_00292_));
 sky130_fd_sc_hd__o21ai_2 _16032_ (.A1(_11255_),
    .A2(latched_store),
    .B1(_10652_),
    .Y(_12053_));
 sky130_fd_sc_hd__o211a_2 _16033_ (.A1(_00292_),
    .A2(_12053_),
    .B1(_11110_),
    .C1(\reg_next_pc[0] ),
    .X(_02770_));
 sky130_fd_sc_hd__and2_2 _16034_ (.A(_11117_),
    .B(_00008_),
    .X(_02769_));
 sky130_fd_sc_hd__and2_2 _16035_ (.A(_11117_),
    .B(_12982_),
    .X(_02768_));
 sky130_fd_sc_hd__buf_1 _16036_ (.A(_11114_),
    .X(_12054_));
 sky130_fd_sc_hd__and2_2 _16037_ (.A(_12054_),
    .B(_00031_),
    .X(_02767_));
 sky130_fd_sc_hd__and2_2 _16038_ (.A(_12054_),
    .B(_00032_),
    .X(_02766_));
 sky130_fd_sc_hd__and2_2 _16039_ (.A(_12054_),
    .B(_00033_),
    .X(_02765_));
 sky130_fd_sc_hd__and2_2 _16040_ (.A(_12054_),
    .B(_00034_),
    .X(_02764_));
 sky130_fd_sc_hd__and2_2 _16041_ (.A(_12054_),
    .B(_00035_),
    .X(_02763_));
 sky130_fd_sc_hd__and2_2 _16042_ (.A(_12054_),
    .B(_00036_),
    .X(_02762_));
 sky130_fd_sc_hd__buf_1 _16043_ (.A(_11114_),
    .X(_12055_));
 sky130_fd_sc_hd__and2_2 _16044_ (.A(_12055_),
    .B(_00037_),
    .X(_02761_));
 sky130_fd_sc_hd__and2_2 _16045_ (.A(_12055_),
    .B(_00009_),
    .X(_02760_));
 sky130_fd_sc_hd__and2_2 _16046_ (.A(_12055_),
    .B(_00010_),
    .X(_02759_));
 sky130_fd_sc_hd__and2_2 _16047_ (.A(_12055_),
    .B(_00011_),
    .X(_02758_));
 sky130_fd_sc_hd__and2_2 _16048_ (.A(_12055_),
    .B(_00012_),
    .X(_02757_));
 sky130_fd_sc_hd__and2_2 _16049_ (.A(_12055_),
    .B(_00013_),
    .X(_02756_));
 sky130_fd_sc_hd__buf_1 _16050_ (.A(_11114_),
    .X(_12056_));
 sky130_fd_sc_hd__and2_2 _16051_ (.A(_12056_),
    .B(_00014_),
    .X(_02755_));
 sky130_fd_sc_hd__and2_2 _16052_ (.A(_12056_),
    .B(_00015_),
    .X(_02754_));
 sky130_fd_sc_hd__and2_2 _16053_ (.A(_12056_),
    .B(_00016_),
    .X(_02753_));
 sky130_fd_sc_hd__and2_2 _16054_ (.A(_12056_),
    .B(_00017_),
    .X(_02752_));
 sky130_fd_sc_hd__and2_2 _16055_ (.A(_12056_),
    .B(_00018_),
    .X(_02751_));
 sky130_fd_sc_hd__and2_2 _16056_ (.A(_12056_),
    .B(_00019_),
    .X(_02750_));
 sky130_fd_sc_hd__buf_1 _16057_ (.A(_10466_),
    .X(_12057_));
 sky130_fd_sc_hd__and2_2 _16058_ (.A(_12057_),
    .B(_00020_),
    .X(_02749_));
 sky130_fd_sc_hd__and2_2 _16059_ (.A(_12057_),
    .B(_00021_),
    .X(_02748_));
 sky130_fd_sc_hd__and2_2 _16060_ (.A(_12057_),
    .B(_00022_),
    .X(_02747_));
 sky130_fd_sc_hd__and2_2 _16061_ (.A(_12057_),
    .B(_00023_),
    .X(_02746_));
 sky130_fd_sc_hd__and2_2 _16062_ (.A(_12057_),
    .B(_00024_),
    .X(_02745_));
 sky130_fd_sc_hd__and2_2 _16063_ (.A(_12057_),
    .B(_00025_),
    .X(_02744_));
 sky130_fd_sc_hd__and2_2 _16064_ (.A(_10464_),
    .B(_00026_),
    .X(_02743_));
 sky130_fd_sc_hd__and2_2 _16065_ (.A(_10464_),
    .B(_00027_),
    .X(_02742_));
 sky130_fd_sc_hd__and2_2 _16066_ (.A(_10464_),
    .B(_00028_),
    .X(_02741_));
 sky130_fd_sc_hd__and2_2 _16067_ (.A(_10464_),
    .B(_00029_),
    .X(_02740_));
 sky130_fd_sc_hd__and2_2 _16068_ (.A(_10464_),
    .B(_00030_),
    .X(_02739_));
 sky130_vsdinv _16069_ (.A(\decoded_imm[1] ),
    .Y(_12058_));
 sky130_vsdinv _16070_ (.A(\mem_rdata_q[8] ),
    .Y(_12059_));
 sky130_fd_sc_hd__nor2_2 _16071_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(_10665_),
    .Y(_12060_));
 sky130_vsdinv _16072_ (.A(\decoded_imm_uj[1] ),
    .Y(_12061_));
 sky130_fd_sc_hd__buf_1 _16073_ (.A(_11793_),
    .X(_12062_));
 sky130_fd_sc_hd__or2_2 _16074_ (.A(_12061_),
    .B(_12062_),
    .X(_12063_));
 sky130_fd_sc_hd__o221a_2 _16075_ (.A1(_12059_),
    .A2(_12060_),
    .B1(_11758_),
    .B2(_11720_),
    .C1(_12063_),
    .X(_12064_));
 sky130_fd_sc_hd__o22ai_2 _16076_ (.A1(_12058_),
    .A2(_11716_),
    .B1(_11701_),
    .B2(_12064_),
    .Y(_02738_));
 sky130_vsdinv _16077_ (.A(\decoded_imm[2] ),
    .Y(_12065_));
 sky130_vsdinv _16078_ (.A(\mem_rdata_q[9] ),
    .Y(_12066_));
 sky130_vsdinv _16079_ (.A(\mem_rdata_q[22] ),
    .Y(_12067_));
 sky130_vsdinv _16080_ (.A(\decoded_imm_uj[2] ),
    .Y(_12068_));
 sky130_fd_sc_hd__or2_2 _16081_ (.A(_12068_),
    .B(_12062_),
    .X(_12069_));
 sky130_fd_sc_hd__o221a_2 _16082_ (.A1(_12066_),
    .A2(_12060_),
    .B1(_12067_),
    .B2(_11720_),
    .C1(_12069_),
    .X(_12070_));
 sky130_fd_sc_hd__o22ai_2 _16083_ (.A1(_12065_),
    .A2(_11716_),
    .B1(_11701_),
    .B2(_12070_),
    .Y(_02737_));
 sky130_vsdinv _16084_ (.A(\decoded_imm[3] ),
    .Y(_12071_));
 sky130_vsdinv _16085_ (.A(\mem_rdata_q[10] ),
    .Y(_12072_));
 sky130_vsdinv _16086_ (.A(\mem_rdata_q[23] ),
    .Y(_12073_));
 sky130_vsdinv _16087_ (.A(\decoded_imm_uj[3] ),
    .Y(_12074_));
 sky130_fd_sc_hd__or2_2 _16088_ (.A(_12074_),
    .B(_12062_),
    .X(_12075_));
 sky130_fd_sc_hd__o221a_2 _16089_ (.A1(_12072_),
    .A2(_12060_),
    .B1(_12073_),
    .B2(_11720_),
    .C1(_12075_),
    .X(_12076_));
 sky130_fd_sc_hd__o22ai_2 _16090_ (.A1(_12071_),
    .A2(_11716_),
    .B1(_11701_),
    .B2(_12076_),
    .Y(_02736_));
 sky130_vsdinv _16091_ (.A(\decoded_imm[4] ),
    .Y(_12077_));
 sky130_fd_sc_hd__buf_1 _16092_ (.A(_11698_),
    .X(_12078_));
 sky130_fd_sc_hd__buf_1 _16093_ (.A(_10760_),
    .X(_12079_));
 sky130_vsdinv _16094_ (.A(\mem_rdata_q[11] ),
    .Y(_12080_));
 sky130_vsdinv _16095_ (.A(\mem_rdata_q[24] ),
    .Y(_12081_));
 sky130_fd_sc_hd__inv_2 _16096_ (.A(\decoded_imm_uj[4] ),
    .Y(_00367_));
 sky130_fd_sc_hd__or2_2 _16097_ (.A(_00367_),
    .B(_12062_),
    .X(_12082_));
 sky130_fd_sc_hd__o221a_2 _16098_ (.A1(_12080_),
    .A2(_12060_),
    .B1(_12081_),
    .B2(_11720_),
    .C1(_12082_),
    .X(_12083_));
 sky130_fd_sc_hd__o22ai_2 _16099_ (.A1(_12077_),
    .A2(_12078_),
    .B1(_12079_),
    .B2(_12083_),
    .Y(_02735_));
 sky130_vsdinv _16100_ (.A(\decoded_imm[5] ),
    .Y(_12084_));
 sky130_vsdinv _16101_ (.A(\decoded_imm_uj[5] ),
    .Y(_12085_));
 sky130_fd_sc_hd__or3_2 _16102_ (.A(is_sb_sh_sw),
    .B(_11719_),
    .C(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_12086_));
 sky130_vsdinv _16103_ (.A(_12086_),
    .Y(_12087_));
 sky130_fd_sc_hd__buf_1 _16104_ (.A(_12087_),
    .X(_12088_));
 sky130_fd_sc_hd__o22a_2 _16105_ (.A1(_12085_),
    .A2(_00323_),
    .B1(_11731_),
    .B2(_12088_),
    .X(_12089_));
 sky130_fd_sc_hd__o22ai_2 _16106_ (.A1(_12084_),
    .A2(_12078_),
    .B1(_12079_),
    .B2(_12089_),
    .Y(_02734_));
 sky130_vsdinv _16107_ (.A(\decoded_imm[6] ),
    .Y(_12090_));
 sky130_fd_sc_hd__buf_1 _16108_ (.A(_12090_),
    .X(_12091_));
 sky130_fd_sc_hd__o2bb2a_2 _16109_ (.A1_N(\decoded_imm_uj[6] ),
    .A2_N(instr_jal),
    .B1(_11739_),
    .B2(_12088_),
    .X(_12092_));
 sky130_fd_sc_hd__o22ai_2 _16110_ (.A1(_12091_),
    .A2(_12078_),
    .B1(_12079_),
    .B2(_12092_),
    .Y(_02733_));
 sky130_vsdinv _16111_ (.A(\decoded_imm[7] ),
    .Y(_12093_));
 sky130_vsdinv _16112_ (.A(\decoded_imm_uj[7] ),
    .Y(_12094_));
 sky130_fd_sc_hd__o22a_2 _16113_ (.A1(_12094_),
    .A2(_00323_),
    .B1(_11723_),
    .B2(_12088_),
    .X(_12095_));
 sky130_fd_sc_hd__o22ai_2 _16114_ (.A1(_12093_),
    .A2(_12078_),
    .B1(_12079_),
    .B2(_12095_),
    .Y(_02732_));
 sky130_vsdinv _16115_ (.A(\decoded_imm[8] ),
    .Y(_12096_));
 sky130_fd_sc_hd__buf_1 _16116_ (.A(_12096_),
    .X(_12097_));
 sky130_vsdinv _16117_ (.A(\decoded_imm_uj[8] ),
    .Y(_12098_));
 sky130_vsdinv _16118_ (.A(_11729_),
    .Y(_12099_));
 sky130_fd_sc_hd__o22a_2 _16119_ (.A1(_12098_),
    .A2(_00323_),
    .B1(_12099_),
    .B2(_12088_),
    .X(_12100_));
 sky130_fd_sc_hd__o22ai_2 _16120_ (.A1(_12097_),
    .A2(_12078_),
    .B1(_12079_),
    .B2(_12100_),
    .Y(_02731_));
 sky130_vsdinv _16121_ (.A(\decoded_imm[9] ),
    .Y(_12101_));
 sky130_vsdinv _16122_ (.A(\decoded_imm_uj[9] ),
    .Y(_12102_));
 sky130_vsdinv _16123_ (.A(_10740_),
    .Y(_12103_));
 sky130_fd_sc_hd__o22a_2 _16124_ (.A1(_12102_),
    .A2(_00323_),
    .B1(_12103_),
    .B2(_12088_),
    .X(_12104_));
 sky130_fd_sc_hd__o22ai_2 _16125_ (.A1(_12101_),
    .A2(_12078_),
    .B1(_12079_),
    .B2(_12104_),
    .Y(_02730_));
 sky130_vsdinv _16126_ (.A(\decoded_imm[10] ),
    .Y(_12105_));
 sky130_fd_sc_hd__buf_1 _16127_ (.A(_11698_),
    .X(_12106_));
 sky130_fd_sc_hd__buf_1 _16128_ (.A(_10760_),
    .X(_12107_));
 sky130_vsdinv _16129_ (.A(\decoded_imm_uj[10] ),
    .Y(_12108_));
 sky130_fd_sc_hd__buf_1 _16130_ (.A(_12062_),
    .X(_12109_));
 sky130_fd_sc_hd__o22a_2 _16131_ (.A1(_12108_),
    .A2(_12109_),
    .B1(_10743_),
    .B2(_12088_),
    .X(_12110_));
 sky130_fd_sc_hd__o22ai_2 _16132_ (.A1(_12105_),
    .A2(_12106_),
    .B1(_12107_),
    .B2(_12110_),
    .Y(_02729_));
 sky130_vsdinv _16133_ (.A(\decoded_imm[11] ),
    .Y(_12111_));
 sky130_vsdinv _16134_ (.A(\decoded_imm_uj[11] ),
    .Y(_12112_));
 sky130_fd_sc_hd__o21ai_2 _16135_ (.A1(_10665_),
    .A2(_11719_),
    .B1(_10742_),
    .Y(_12113_));
 sky130_fd_sc_hd__o221a_2 _16136_ (.A1(_12112_),
    .A2(_12109_),
    .B1(_10607_),
    .B2(_11717_),
    .C1(_12113_),
    .X(_12114_));
 sky130_fd_sc_hd__o22ai_2 _16137_ (.A1(_12111_),
    .A2(_12106_),
    .B1(_12107_),
    .B2(_12114_),
    .Y(_02728_));
 sky130_vsdinv _16138_ (.A(\decoded_imm[12] ),
    .Y(_12115_));
 sky130_vsdinv _16139_ (.A(\decoded_imm_uj[12] ),
    .Y(_12116_));
 sky130_vsdinv _16140_ (.A(_10630_),
    .Y(_12117_));
 sky130_fd_sc_hd__buf_1 _16141_ (.A(_12117_),
    .X(_12118_));
 sky130_fd_sc_hd__or2_2 _16142_ (.A(_11761_),
    .B(_12087_),
    .X(_12119_));
 sky130_fd_sc_hd__buf_1 _16143_ (.A(_12119_),
    .X(_12120_));
 sky130_fd_sc_hd__o221a_2 _16144_ (.A1(_12116_),
    .A2(_12109_),
    .B1(_10726_),
    .B2(_12118_),
    .C1(_12120_),
    .X(_12121_));
 sky130_fd_sc_hd__o22ai_2 _16145_ (.A1(_12115_),
    .A2(_12106_),
    .B1(_12107_),
    .B2(_12121_),
    .Y(_02727_));
 sky130_vsdinv _16146_ (.A(\decoded_imm[13] ),
    .Y(_12122_));
 sky130_vsdinv _16147_ (.A(\decoded_imm_uj[13] ),
    .Y(_12123_));
 sky130_fd_sc_hd__buf_1 _16148_ (.A(_12117_),
    .X(_12124_));
 sky130_fd_sc_hd__o221a_2 _16149_ (.A1(_12123_),
    .A2(_12109_),
    .B1(_10724_),
    .B2(_12124_),
    .C1(_12120_),
    .X(_12125_));
 sky130_fd_sc_hd__o22ai_2 _16150_ (.A1(_12122_),
    .A2(_12106_),
    .B1(_12107_),
    .B2(_12125_),
    .Y(_02726_));
 sky130_vsdinv _16151_ (.A(\decoded_imm[14] ),
    .Y(_12126_));
 sky130_vsdinv _16152_ (.A(\decoded_imm_uj[14] ),
    .Y(_12127_));
 sky130_fd_sc_hd__o221a_2 _16153_ (.A1(_12127_),
    .A2(_12109_),
    .B1(_00334_),
    .B2(_12124_),
    .C1(_12120_),
    .X(_12128_));
 sky130_fd_sc_hd__o22ai_2 _16154_ (.A1(_12126_),
    .A2(_12106_),
    .B1(_12107_),
    .B2(_12128_),
    .Y(_02725_));
 sky130_vsdinv _16155_ (.A(\decoded_imm[15] ),
    .Y(_12129_));
 sky130_vsdinv _16156_ (.A(\decoded_imm_uj[15] ),
    .Y(_12130_));
 sky130_vsdinv _16157_ (.A(\mem_rdata_q[15] ),
    .Y(_12131_));
 sky130_fd_sc_hd__o221a_2 _16158_ (.A1(_12130_),
    .A2(_11794_),
    .B1(_12131_),
    .B2(_12124_),
    .C1(_12120_),
    .X(_12132_));
 sky130_fd_sc_hd__o22ai_2 _16159_ (.A1(_12129_),
    .A2(_12106_),
    .B1(_12107_),
    .B2(_12132_),
    .Y(_02724_));
 sky130_vsdinv _16160_ (.A(\decoded_imm[16] ),
    .Y(_12133_));
 sky130_fd_sc_hd__buf_1 _16161_ (.A(_12133_),
    .X(_12134_));
 sky130_vsdinv _16162_ (.A(\decoded_imm_uj[16] ),
    .Y(_12135_));
 sky130_vsdinv _16163_ (.A(\mem_rdata_q[16] ),
    .Y(_12136_));
 sky130_fd_sc_hd__o221a_2 _16164_ (.A1(_12135_),
    .A2(_11794_),
    .B1(_12136_),
    .B2(_12124_),
    .C1(_12120_),
    .X(_12137_));
 sky130_fd_sc_hd__o22ai_2 _16165_ (.A1(_12134_),
    .A2(_11798_),
    .B1(_11107_),
    .B2(_12137_),
    .Y(_02723_));
 sky130_vsdinv _16166_ (.A(\decoded_imm[17] ),
    .Y(_12138_));
 sky130_vsdinv _16167_ (.A(\decoded_imm_uj[17] ),
    .Y(_12139_));
 sky130_vsdinv _16168_ (.A(\mem_rdata_q[17] ),
    .Y(_12140_));
 sky130_fd_sc_hd__o221a_2 _16169_ (.A1(_12139_),
    .A2(_11794_),
    .B1(_12140_),
    .B2(_12124_),
    .C1(_12120_),
    .X(_12141_));
 sky130_fd_sc_hd__o22ai_2 _16170_ (.A1(_12138_),
    .A2(_11798_),
    .B1(_11107_),
    .B2(_12141_),
    .Y(_02722_));
 sky130_vsdinv _16171_ (.A(\decoded_imm[18] ),
    .Y(_12142_));
 sky130_vsdinv _16172_ (.A(\decoded_imm_uj[18] ),
    .Y(_12143_));
 sky130_vsdinv _16173_ (.A(\mem_rdata_q[18] ),
    .Y(_12144_));
 sky130_fd_sc_hd__o221a_2 _16174_ (.A1(_12143_),
    .A2(_11794_),
    .B1(_12144_),
    .B2(_12124_),
    .C1(_12119_),
    .X(_12145_));
 sky130_fd_sc_hd__o22ai_2 _16175_ (.A1(_12142_),
    .A2(_11798_),
    .B1(_11107_),
    .B2(_12145_),
    .Y(_02721_));
 sky130_vsdinv _16176_ (.A(\decoded_imm[19] ),
    .Y(_12146_));
 sky130_vsdinv _16177_ (.A(\decoded_imm_uj[19] ),
    .Y(_12147_));
 sky130_vsdinv _16178_ (.A(\mem_rdata_q[19] ),
    .Y(_12148_));
 sky130_fd_sc_hd__o221a_2 _16179_ (.A1(_12147_),
    .A2(_11794_),
    .B1(_12148_),
    .B2(_12117_),
    .C1(_12119_),
    .X(_12149_));
 sky130_fd_sc_hd__o22ai_2 _16180_ (.A1(_12146_),
    .A2(_11798_),
    .B1(_11107_),
    .B2(_12149_),
    .Y(_02720_));
 sky130_fd_sc_hd__nor2_2 _16181_ (.A(_11761_),
    .B(_11720_),
    .Y(_12150_));
 sky130_fd_sc_hd__buf_1 _16182_ (.A(_12150_),
    .X(_12151_));
 sky130_fd_sc_hd__buf_1 _16183_ (.A(_12117_),
    .X(_12152_));
 sky130_fd_sc_hd__o21ai_2 _16184_ (.A1(_11718_),
    .A2(_12152_),
    .B1(_11788_),
    .Y(_12153_));
 sky130_vsdinv _16185_ (.A(\decoded_imm_uj[20] ),
    .Y(_12154_));
 sky130_fd_sc_hd__buf_1 _16186_ (.A(_12154_),
    .X(_12155_));
 sky130_fd_sc_hd__buf_1 _16187_ (.A(_12155_),
    .X(_12156_));
 sky130_fd_sc_hd__buf_1 _16188_ (.A(_12156_),
    .X(_12157_));
 sky130_fd_sc_hd__buf_1 _16189_ (.A(_12157_),
    .X(_12158_));
 sky130_fd_sc_hd__o22ai_2 _16190_ (.A1(_12158_),
    .A2(_12062_),
    .B1(_11761_),
    .B2(_12060_),
    .Y(_12159_));
 sky130_fd_sc_hd__buf_1 _16191_ (.A(_12159_),
    .X(_12160_));
 sky130_fd_sc_hd__o32a_2 _16192_ (.A1(_12151_),
    .A2(_12153_),
    .A3(_12160_),
    .B1(\decoded_imm[20] ),
    .B2(_11699_),
    .X(_02719_));
 sky130_fd_sc_hd__o21ai_2 _16193_ (.A1(_11758_),
    .A2(_12152_),
    .B1(_11788_),
    .Y(_12161_));
 sky130_fd_sc_hd__o32a_2 _16194_ (.A1(_12151_),
    .A2(_12161_),
    .A3(_12160_),
    .B1(\decoded_imm[21] ),
    .B2(_11699_),
    .X(_02718_));
 sky130_fd_sc_hd__o21ai_2 _16195_ (.A1(_12067_),
    .A2(_12152_),
    .B1(_11788_),
    .Y(_12162_));
 sky130_fd_sc_hd__o32a_2 _16196_ (.A1(_12151_),
    .A2(_12162_),
    .A3(_12160_),
    .B1(\decoded_imm[22] ),
    .B2(_11699_),
    .X(_02717_));
 sky130_fd_sc_hd__o21ai_2 _16197_ (.A1(_12073_),
    .A2(_12152_),
    .B1(_11788_),
    .Y(_12163_));
 sky130_fd_sc_hd__o32a_2 _16198_ (.A1(_12151_),
    .A2(_12163_),
    .A3(_12160_),
    .B1(\decoded_imm[23] ),
    .B2(_11699_),
    .X(_02716_));
 sky130_fd_sc_hd__buf_1 _16199_ (.A(_10748_),
    .X(_12164_));
 sky130_fd_sc_hd__o21ai_2 _16200_ (.A1(_12081_),
    .A2(_12152_),
    .B1(_12164_),
    .Y(_12165_));
 sky130_fd_sc_hd__o32a_2 _16201_ (.A1(_12151_),
    .A2(_12165_),
    .A3(_12160_),
    .B1(\decoded_imm[24] ),
    .B2(_11699_),
    .X(_02715_));
 sky130_fd_sc_hd__o21ai_2 _16202_ (.A1(_11731_),
    .A2(_12152_),
    .B1(_12164_),
    .Y(_12166_));
 sky130_fd_sc_hd__buf_1 _16203_ (.A(_11698_),
    .X(_12167_));
 sky130_fd_sc_hd__o32a_2 _16204_ (.A1(_12151_),
    .A2(_12166_),
    .A3(_12160_),
    .B1(\decoded_imm[25] ),
    .B2(_12167_),
    .X(_02714_));
 sky130_fd_sc_hd__o21ai_2 _16205_ (.A1(_11739_),
    .A2(_12118_),
    .B1(_12164_),
    .Y(_12168_));
 sky130_fd_sc_hd__o32a_2 _16206_ (.A1(_12150_),
    .A2(_12168_),
    .A3(_12159_),
    .B1(\decoded_imm[26] ),
    .B2(_12167_),
    .X(_02713_));
 sky130_fd_sc_hd__o21ai_2 _16207_ (.A1(_11723_),
    .A2(_12118_),
    .B1(_12164_),
    .Y(_12169_));
 sky130_fd_sc_hd__o32a_2 _16208_ (.A1(_12150_),
    .A2(_12169_),
    .A3(_12159_),
    .B1(\decoded_imm[27] ),
    .B2(_12167_),
    .X(_02712_));
 sky130_fd_sc_hd__o21ai_2 _16209_ (.A1(_12099_),
    .A2(_12118_),
    .B1(_12164_),
    .Y(_12170_));
 sky130_fd_sc_hd__o32a_2 _16210_ (.A1(_12150_),
    .A2(_12170_),
    .A3(_12159_),
    .B1(\decoded_imm[28] ),
    .B2(_12167_),
    .X(_02711_));
 sky130_fd_sc_hd__o21ai_2 _16211_ (.A1(_12103_),
    .A2(_12118_),
    .B1(_12164_),
    .Y(_12171_));
 sky130_fd_sc_hd__o32a_2 _16212_ (.A1(_12150_),
    .A2(_12171_),
    .A3(_12159_),
    .B1(\decoded_imm[29] ),
    .B2(_12167_),
    .X(_02710_));
 sky130_fd_sc_hd__o21ai_2 _16213_ (.A1(_10743_),
    .A2(_12118_),
    .B1(_10749_),
    .Y(_12172_));
 sky130_fd_sc_hd__o32a_2 _16214_ (.A1(_12150_),
    .A2(_12172_),
    .A3(_12159_),
    .B1(\decoded_imm[30] ),
    .B2(_12167_),
    .X(_02709_));
 sky130_vsdinv _16215_ (.A(\decoded_imm[31] ),
    .Y(_12173_));
 sky130_fd_sc_hd__buf_1 _16216_ (.A(_12158_),
    .X(_12174_));
 sky130_fd_sc_hd__nor2_2 _16217_ (.A(_10630_),
    .B(_12086_),
    .Y(_12175_));
 sky130_fd_sc_hd__o22a_2 _16218_ (.A1(_12174_),
    .A2(_12109_),
    .B1(_11761_),
    .B2(_12175_),
    .X(_12176_));
 sky130_fd_sc_hd__o22ai_2 _16219_ (.A1(_12173_),
    .A2(_11798_),
    .B1(_11107_),
    .B2(_12176_),
    .Y(_02708_));
 sky130_fd_sc_hd__or2_2 _16220_ (.A(\cpu_state[4] ),
    .B(\cpu_state[2] ),
    .X(_12177_));
 sky130_fd_sc_hd__buf_1 _16221_ (.A(_12177_),
    .X(_02542_));
 sky130_vsdinv _16222_ (.A(_02542_),
    .Y(_12178_));
 sky130_fd_sc_hd__or4_2 _16223_ (.A(_10477_),
    .B(_00331_),
    .C(_11426_),
    .D(_10614_),
    .X(_12179_));
 sky130_vsdinv _16224_ (.A(_12179_),
    .Y(_12180_));
 sky130_fd_sc_hd__a32o_2 _16225_ (.A1(_12942_),
    .A2(_12178_),
    .A3(_12180_),
    .B1(\latched_rd[0] ),
    .B2(_12179_),
    .X(_02707_));
 sky130_fd_sc_hd__nor2_2 _16226_ (.A(_00308_),
    .B(_02542_),
    .Y(_12181_));
 sky130_fd_sc_hd__a32o_2 _16227_ (.A1(\decoded_rd[1] ),
    .A2(_12180_),
    .A3(_12181_),
    .B1(\latched_rd[1] ),
    .B2(_12179_),
    .X(_02706_));
 sky130_fd_sc_hd__a32o_2 _16228_ (.A1(\decoded_rd[2] ),
    .A2(_12180_),
    .A3(_12181_),
    .B1(_11310_),
    .B2(_12179_),
    .X(_02705_));
 sky130_fd_sc_hd__a32o_2 _16229_ (.A1(\decoded_rd[3] ),
    .A2(_12180_),
    .A3(_12181_),
    .B1(_11252_),
    .B2(_12179_),
    .X(_02704_));
 sky130_fd_sc_hd__buf_1 _16230_ (.A(_11082_),
    .X(_12182_));
 sky130_fd_sc_hd__or3_2 _16231_ (.A(_10665_),
    .B(_12182_),
    .C(_00310_),
    .X(_12183_));
 sky130_fd_sc_hd__o31ai_2 _16232_ (.A1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2(is_slli_srli_srai),
    .A3(is_lui_auipc_jal),
    .B1(_10614_),
    .Y(_12184_));
 sky130_fd_sc_hd__a21oi_2 _16233_ (.A1(_12183_),
    .A2(_12184_),
    .B1(_11330_),
    .Y(_02703_));
 sky130_vsdinv _16234_ (.A(mem_la_wdata[4]),
    .Y(_12185_));
 sky130_fd_sc_hd__buf_1 _16235_ (.A(_12185_),
    .X(_02327_));
 sky130_fd_sc_hd__and2_2 _16236_ (.A(_02327_),
    .B(_02558_),
    .X(_02702_));
 sky130_fd_sc_hd__and2_2 _16237_ (.A(_02327_),
    .B(_02557_),
    .X(_02701_));
 sky130_fd_sc_hd__and2_2 _16238_ (.A(_02327_),
    .B(_02556_),
    .X(_02700_));
 sky130_fd_sc_hd__buf_1 _16239_ (.A(_12185_),
    .X(_12186_));
 sky130_fd_sc_hd__and2_2 _16240_ (.A(_12186_),
    .B(_02555_),
    .X(_02699_));
 sky130_fd_sc_hd__and2_2 _16241_ (.A(_12186_),
    .B(_02554_),
    .X(_02698_));
 sky130_fd_sc_hd__and2_2 _16242_ (.A(_12186_),
    .B(_02553_),
    .X(_02697_));
 sky130_fd_sc_hd__and2_2 _16243_ (.A(_12186_),
    .B(_02552_),
    .X(_02696_));
 sky130_fd_sc_hd__and2_2 _16244_ (.A(_12186_),
    .B(_02551_),
    .X(_02695_));
 sky130_vsdinv _16245_ (.A(mem_la_wdata[3]),
    .Y(_12187_));
 sky130_fd_sc_hd__buf_1 _16246_ (.A(_12187_),
    .X(_12188_));
 sky130_fd_sc_hd__buf_1 _16247_ (.A(_12188_),
    .X(_02324_));
 sky130_fd_sc_hd__and2_2 _16248_ (.A(_02324_),
    .B(_00122_),
    .X(_02550_));
 sky130_fd_sc_hd__buf_1 _16249_ (.A(_12187_),
    .X(_12189_));
 sky130_fd_sc_hd__and3_2 _16250_ (.A(_12189_),
    .B(_00122_),
    .C(_12186_),
    .X(_02694_));
 sky130_fd_sc_hd__and2_2 _16251_ (.A(_02324_),
    .B(_00116_),
    .X(_02549_));
 sky130_fd_sc_hd__buf_1 _16252_ (.A(_12185_),
    .X(_12190_));
 sky130_fd_sc_hd__and3_2 _16253_ (.A(_12189_),
    .B(_00116_),
    .C(_12190_),
    .X(_02693_));
 sky130_fd_sc_hd__and2_2 _16254_ (.A(_02324_),
    .B(_00110_),
    .X(_02548_));
 sky130_fd_sc_hd__and3_2 _16255_ (.A(_12189_),
    .B(_00110_),
    .C(_12190_),
    .X(_02692_));
 sky130_fd_sc_hd__and2_2 _16256_ (.A(_02324_),
    .B(_00104_),
    .X(_02547_));
 sky130_fd_sc_hd__and3_2 _16257_ (.A(_12189_),
    .B(_00104_),
    .C(_12190_),
    .X(_02691_));
 sky130_vsdinv _16258_ (.A(mem_la_wdata[2]),
    .Y(_12191_));
 sky130_fd_sc_hd__buf_1 _16259_ (.A(_12191_),
    .X(_02321_));
 sky130_fd_sc_hd__and3_2 _16260_ (.A(_02321_),
    .B(_00094_),
    .C(_12188_),
    .X(_02546_));
 sky130_fd_sc_hd__and2_2 _16261_ (.A(_02321_),
    .B(_00094_),
    .X(_00095_));
 sky130_fd_sc_hd__and3_2 _16262_ (.A(_12189_),
    .B(_00095_),
    .C(_12190_),
    .X(_02690_));
 sky130_fd_sc_hd__and3_2 _16263_ (.A(_02321_),
    .B(_00084_),
    .C(_12188_),
    .X(_02545_));
 sky130_fd_sc_hd__and2_2 _16264_ (.A(_12191_),
    .B(_00084_),
    .X(_00085_));
 sky130_fd_sc_hd__and3_2 _16265_ (.A(_12189_),
    .B(_00085_),
    .C(_12190_),
    .X(_02689_));
 sky130_vsdinv _16266_ (.A(mem_la_wdata[1]),
    .Y(_12192_));
 sky130_fd_sc_hd__buf_1 _16267_ (.A(_12192_),
    .X(_02318_));
 sky130_fd_sc_hd__and3_2 _16268_ (.A(_02318_),
    .B(_00066_),
    .C(_12191_),
    .X(_12193_));
 sky130_fd_sc_hd__buf_1 _16269_ (.A(_12193_),
    .X(_00068_));
 sky130_fd_sc_hd__nand2_2 _16270_ (.A(_12188_),
    .B(_00068_),
    .Y(_12194_));
 sky130_vsdinv _16271_ (.A(_12194_),
    .Y(_02544_));
 sky130_fd_sc_hd__nor2_2 _16272_ (.A(_11360_),
    .B(_12194_),
    .Y(_02688_));
 sky130_vsdinv _16273_ (.A(pcpi_rs1[0]),
    .Y(_12195_));
 sky130_fd_sc_hd__buf_1 _16274_ (.A(_12195_),
    .X(_12196_));
 sky130_fd_sc_hd__nor2_2 _16275_ (.A(_11364_),
    .B(_12196_),
    .Y(_00048_));
 sky130_fd_sc_hd__nand2_2 _16276_ (.A(_12192_),
    .B(_00048_),
    .Y(_12197_));
 sky130_fd_sc_hd__inv_2 _16277_ (.A(_12197_),
    .Y(_00049_));
 sky130_fd_sc_hd__and3_2 _16278_ (.A(_02321_),
    .B(_00049_),
    .C(_12188_),
    .X(_02543_));
 sky130_fd_sc_hd__nor2_2 _16279_ (.A(_11362_),
    .B(_12197_),
    .Y(_00050_));
 sky130_fd_sc_hd__and3_2 _16280_ (.A(_12188_),
    .B(_00050_),
    .C(_12190_),
    .X(_02687_));
 sky130_fd_sc_hd__o211a_2 _16281_ (.A1(\reg_pc[1] ),
    .A2(\reg_next_pc[0] ),
    .B1(resetn),
    .C1(mem_do_rinst),
    .X(_12198_));
 sky130_fd_sc_hd__buf_1 _16282_ (.A(_12198_),
    .X(_00307_));
 sky130_fd_sc_hd__or2_2 _16283_ (.A(irq_active),
    .B(\irq_mask[2] ),
    .X(_12199_));
 sky130_fd_sc_hd__buf_1 _16284_ (.A(_12199_),
    .X(_12200_));
 sky130_fd_sc_hd__buf_1 _16285_ (.A(_12200_),
    .X(_12201_));
 sky130_fd_sc_hd__nor2_2 _16286_ (.A(_11111_),
    .B(_12201_),
    .Y(_00312_));
 sky130_fd_sc_hd__o21ai_2 _16287_ (.A1(mem_do_wdata),
    .A2(mem_do_rdata),
    .B1(resetn),
    .Y(_12202_));
 sky130_fd_sc_hd__inv_2 _16288_ (.A(_12202_),
    .Y(_00303_));
 sky130_vsdinv _16289_ (.A(_12198_),
    .Y(_12203_));
 sky130_fd_sc_hd__or2_2 _16290_ (.A(_12203_),
    .B(_12199_),
    .X(_12204_));
 sky130_fd_sc_hd__o21a_2 _16291_ (.A1(decoder_trigger),
    .A2(_11103_),
    .B1(_10564_),
    .X(_12205_));
 sky130_fd_sc_hd__buf_1 _16292_ (.A(_12202_),
    .X(_12206_));
 sky130_vsdinv _16293_ (.A(\mem_wordsize[2] ),
    .Y(_12207_));
 sky130_fd_sc_hd__or2_2 _16294_ (.A(_12196_),
    .B(_12207_),
    .X(_12208_));
 sky130_fd_sc_hd__inv_2 _16295_ (.A(_12208_),
    .Y(_00306_));
 sky130_vsdinv _16296_ (.A(\mem_wordsize[0] ),
    .Y(_12209_));
 sky130_fd_sc_hd__nor2_2 _16297_ (.A(_11861_),
    .B(_11863_),
    .Y(_00304_));
 sky130_fd_sc_hd__or2_2 _16298_ (.A(_12209_),
    .B(_00304_),
    .X(_12210_));
 sky130_fd_sc_hd__or3_2 _16299_ (.A(_11793_),
    .B(_10509_),
    .C(_10565_),
    .X(_12211_));
 sky130_fd_sc_hd__or2_2 _16300_ (.A(_10475_),
    .B(_12211_),
    .X(_12212_));
 sky130_fd_sc_hd__or3_2 _16301_ (.A(decoder_trigger),
    .B(_00309_),
    .C(_11103_),
    .X(_12213_));
 sky130_fd_sc_hd__inv_2 _16302_ (.A(_12210_),
    .Y(_00305_));
 sky130_fd_sc_hd__o32a_2 _16303_ (.A1(_12200_),
    .A2(_12210_),
    .A3(_12212_),
    .B1(_12213_),
    .B2(_00305_),
    .X(_12214_));
 sky130_fd_sc_hd__o41a_2 _16304_ (.A1(_12199_),
    .A2(_12210_),
    .A3(_12206_),
    .A4(_00306_),
    .B1(_00303_),
    .X(_12215_));
 sky130_fd_sc_hd__or2_2 _16305_ (.A(_12213_),
    .B(_12215_),
    .X(_12216_));
 sky130_fd_sc_hd__nor2_2 _16306_ (.A(_00306_),
    .B(_00305_),
    .Y(_12217_));
 sky130_fd_sc_hd__a21oi_2 _16307_ (.A1(_10708_),
    .A2(_10456_),
    .B1(_12217_),
    .Y(_12218_));
 sky130_fd_sc_hd__nand2_2 _16308_ (.A(resetn),
    .B(_00308_),
    .Y(_12219_));
 sky130_fd_sc_hd__or3b_2 _16309_ (.A(_12200_),
    .B(_12219_),
    .C_N(_12218_),
    .X(_12220_));
 sky130_fd_sc_hd__o221a_2 _16310_ (.A1(_11104_),
    .A2(_00303_),
    .B1(_12218_),
    .B2(_12212_),
    .C1(_12220_),
    .X(_12221_));
 sky130_fd_sc_hd__o311a_2 _16311_ (.A1(_12206_),
    .A2(_00306_),
    .A3(_12214_),
    .B1(_12216_),
    .C1(_12221_),
    .X(_12222_));
 sky130_vsdinv _16312_ (.A(_12204_),
    .Y(_12223_));
 sky130_fd_sc_hd__o21a_2 _16313_ (.A1(_12202_),
    .A2(_12217_),
    .B1(_12203_),
    .X(_12224_));
 sky130_fd_sc_hd__nor2_2 _16314_ (.A(_12223_),
    .B(_12224_),
    .Y(_12225_));
 sky130_vsdinv _16315_ (.A(_12199_),
    .Y(_12226_));
 sky130_fd_sc_hd__a31o_2 _16316_ (.A1(_12226_),
    .A2(_00306_),
    .A3(_00303_),
    .B1(_12223_),
    .X(_12227_));
 sky130_vsdinv _16317_ (.A(_12227_),
    .Y(_12228_));
 sky130_fd_sc_hd__or2_2 _16318_ (.A(_12198_),
    .B(_00306_),
    .X(_12229_));
 sky130_fd_sc_hd__or2_2 _16319_ (.A(_12206_),
    .B(_12229_),
    .X(_12230_));
 sky130_fd_sc_hd__a211o_2 _16320_ (.A1(_12201_),
    .A2(_00305_),
    .B1(_12230_),
    .C1(_11104_),
    .X(_12231_));
 sky130_fd_sc_hd__o221a_2 _16321_ (.A1(_12219_),
    .A2(_12225_),
    .B1(_12212_),
    .B2(_12228_),
    .C1(_12231_),
    .X(_12232_));
 sky130_fd_sc_hd__o221a_2 _16322_ (.A1(_12204_),
    .A2(_12205_),
    .B1(_00307_),
    .B2(_12222_),
    .C1(_12232_),
    .X(_12233_));
 sky130_fd_sc_hd__or2_2 _16323_ (.A(_12226_),
    .B(_12224_),
    .X(_12234_));
 sky130_vsdinv _16324_ (.A(_12234_),
    .Y(_12235_));
 sky130_fd_sc_hd__buf_1 _16325_ (.A(_12235_),
    .X(_12236_));
 sky130_fd_sc_hd__or4_2 _16326_ (.A(irq_active),
    .B(\irq_mask[1] ),
    .C(\pcpi_mul.active[1] ),
    .D(_00311_),
    .X(_12237_));
 sky130_fd_sc_hd__o31a_2 _16327_ (.A1(_12200_),
    .A2(_12210_),
    .A3(_12230_),
    .B1(_12225_),
    .X(_12238_));
 sky130_fd_sc_hd__o22a_2 _16328_ (.A1(_10623_),
    .A2(_12236_),
    .B1(_12237_),
    .B2(_12238_),
    .X(_12239_));
 sky130_fd_sc_hd__o21ai_2 _16329_ (.A1(_12226_),
    .A2(_12217_),
    .B1(_12203_),
    .Y(_12240_));
 sky130_fd_sc_hd__or3_2 _16330_ (.A(_12200_),
    .B(_12208_),
    .C(_00307_),
    .X(_12241_));
 sky130_fd_sc_hd__o32a_2 _16331_ (.A1(_10477_),
    .A2(_11083_),
    .A3(_12237_),
    .B1(_10646_),
    .B2(_12213_),
    .X(_12242_));
 sky130_fd_sc_hd__or3_2 _16332_ (.A(_10646_),
    .B(_11104_),
    .C(_12241_),
    .X(_12243_));
 sky130_fd_sc_hd__o221a_2 _16333_ (.A1(_11109_),
    .A2(_12240_),
    .B1(_12241_),
    .B2(_12242_),
    .C1(_12243_),
    .X(_12244_));
 sky130_fd_sc_hd__o21ai_2 _16334_ (.A1(_00307_),
    .A2(_12218_),
    .B1(_12200_),
    .Y(_12245_));
 sky130_fd_sc_hd__nand2_2 _16335_ (.A(_10443_),
    .B(_12245_),
    .Y(_12246_));
 sky130_fd_sc_hd__or4_2 _16336_ (.A(_10606_),
    .B(alu_wait),
    .C(_10609_),
    .D(_10454_),
    .X(_12247_));
 sky130_fd_sc_hd__o21a_2 _16337_ (.A1(_00307_),
    .A2(_00303_),
    .B1(_12204_),
    .X(_12248_));
 sky130_fd_sc_hd__a211oi_2 _16338_ (.A1(_11426_),
    .A2(_12234_),
    .B1(_10477_),
    .C1(_00314_),
    .Y(_12249_));
 sky130_fd_sc_hd__o221a_2 _16339_ (.A1(_12235_),
    .A2(_12247_),
    .B1(_11109_),
    .B2(_12248_),
    .C1(_12249_),
    .X(_12250_));
 sky130_fd_sc_hd__o31a_2 _16340_ (.A1(_11030_),
    .A2(_10621_),
    .A3(_12246_),
    .B1(_12250_),
    .X(_12251_));
 sky130_fd_sc_hd__o221a_2 _16341_ (.A1(_11083_),
    .A2(_12239_),
    .B1(_12206_),
    .B2(_12244_),
    .C1(_12251_),
    .X(_12252_));
 sky130_fd_sc_hd__o21ai_2 _16342_ (.A1(_00322_),
    .A2(_12233_),
    .B1(_12252_),
    .Y(_00039_));
 sky130_fd_sc_hd__nor2_2 _16343_ (.A(_10675_),
    .B(_12246_),
    .Y(_00040_));
 sky130_fd_sc_hd__and3_2 _16344_ (.A(_10457_),
    .B(_12224_),
    .C(_10808_),
    .X(_12253_));
 sky130_fd_sc_hd__a31oi_2 _16345_ (.A1(_11027_),
    .A2(_12234_),
    .A3(_10664_),
    .B1(_12253_),
    .Y(_12254_));
 sky130_fd_sc_hd__buf_1 _16346_ (.A(_10459_),
    .X(_12255_));
 sky130_fd_sc_hd__buf_1 _16347_ (.A(_12255_),
    .X(_12256_));
 sky130_vsdinv _16348_ (.A(mem_do_prefetch),
    .Y(_12257_));
 sky130_fd_sc_hd__or2_2 _16349_ (.A(_12257_),
    .B(_10661_),
    .X(_12258_));
 sky130_fd_sc_hd__or2_2 _16350_ (.A(_10476_),
    .B(_10808_),
    .X(_12259_));
 sky130_vsdinv _16351_ (.A(_11108_),
    .Y(_12260_));
 sky130_fd_sc_hd__or2_2 _16352_ (.A(_12259_),
    .B(_12260_),
    .X(_12261_));
 sky130_fd_sc_hd__o32a_2 _16353_ (.A1(_12201_),
    .A2(_12224_),
    .A3(_12258_),
    .B1(_12236_),
    .B2(_12261_),
    .X(_12262_));
 sky130_fd_sc_hd__o22ai_2 _16354_ (.A1(_10689_),
    .A2(_12254_),
    .B1(_12256_),
    .B2(_12262_),
    .Y(_00044_));
 sky130_fd_sc_hd__nor2_2 _16355_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B(is_slli_srli_srai),
    .Y(_01304_));
 sky130_fd_sc_hd__or4b_2 _16356_ (.A(is_lui_auipc_jal),
    .B(_12235_),
    .C(_10622_),
    .D_N(_01304_),
    .X(_12263_));
 sky130_fd_sc_hd__o32a_2 _16357_ (.A1(_11083_),
    .A2(_11086_),
    .A3(_12236_),
    .B1(_10664_),
    .B2(_12263_),
    .X(_12264_));
 sky130_fd_sc_hd__nor2_2 _16358_ (.A(_11017_),
    .B(_12264_),
    .Y(_00041_));
 sky130_fd_sc_hd__a211o_2 _16359_ (.A1(_10560_),
    .A2(_10510_),
    .B1(\pcpi_mul.active[1] ),
    .C1(_00311_),
    .X(_12265_));
 sky130_fd_sc_hd__or3_2 _16360_ (.A(_11083_),
    .B(_12265_),
    .C(_12236_),
    .X(_12266_));
 sky130_fd_sc_hd__a31oi_2 _16361_ (.A1(_11251_),
    .A2(_12245_),
    .A3(_12266_),
    .B1(_10974_),
    .Y(_00038_));
 sky130_vsdinv _16362_ (.A(_11020_),
    .Y(_00315_));
 sky130_fd_sc_hd__or3_2 _16363_ (.A(_10476_),
    .B(_10666_),
    .C(_12182_),
    .X(_12267_));
 sky130_fd_sc_hd__or3_2 _16364_ (.A(_12206_),
    .B(_12210_),
    .C(_11807_),
    .X(_12268_));
 sky130_fd_sc_hd__o32a_2 _16365_ (.A1(_12201_),
    .A2(_12206_),
    .A3(_12267_),
    .B1(_12258_),
    .B2(_12268_),
    .X(_12269_));
 sky130_fd_sc_hd__o21bai_2 _16366_ (.A1(_12227_),
    .A2(_12224_),
    .B1_N(_12267_),
    .Y(_12270_));
 sky130_fd_sc_hd__a41o_2 _16367_ (.A1(_00303_),
    .A2(_00305_),
    .A3(_12203_),
    .A4(_12208_),
    .B1(_12258_),
    .X(_12271_));
 sky130_fd_sc_hd__a211o_2 _16368_ (.A1(_12261_),
    .A2(_12271_),
    .B1(_11807_),
    .C1(_12236_),
    .X(_12272_));
 sky130_fd_sc_hd__o311a_2 _16369_ (.A1(_12201_),
    .A2(_12229_),
    .A3(_12269_),
    .B1(_12270_),
    .C1(_12272_),
    .X(_12273_));
 sky130_vsdinv _16370_ (.A(_12273_),
    .Y(_00043_));
 sky130_fd_sc_hd__and3_2 _16371_ (.A(_11106_),
    .B(_00290_),
    .C(_10484_),
    .X(mem_la_read));
 sky130_vsdinv _16372_ (.A(_11396_),
    .Y(mem_la_write));
 sky130_fd_sc_hd__nor2_2 _16373_ (.A(_00291_),
    .B(_11807_),
    .Y(_00317_));
 sky130_fd_sc_hd__buf_1 _16374_ (.A(_10610_),
    .X(_12274_));
 sky130_fd_sc_hd__or3_2 _16375_ (.A(_10607_),
    .B(alu_wait),
    .C(_10661_),
    .X(_12275_));
 sky130_fd_sc_hd__o21a_2 _16376_ (.A1(_00305_),
    .A2(_12230_),
    .B1(_12228_),
    .X(_12276_));
 sky130_fd_sc_hd__o32a_2 _16377_ (.A1(_10482_),
    .A2(_00302_),
    .A3(_12236_),
    .B1(_12275_),
    .B2(_12276_),
    .X(_12277_));
 sky130_fd_sc_hd__or2_2 _16378_ (.A(_10609_),
    .B(_12215_),
    .X(_12278_));
 sky130_fd_sc_hd__o32a_2 _16379_ (.A1(_10482_),
    .A2(_12218_),
    .A3(_12183_),
    .B1(_12275_),
    .B2(_12278_),
    .X(_12279_));
 sky130_fd_sc_hd__o32a_2 _16380_ (.A1(_12201_),
    .A2(_12224_),
    .A3(_12183_),
    .B1(_12184_),
    .B2(_12246_),
    .X(_12280_));
 sky130_fd_sc_hd__o221ai_2 _16381_ (.A1(_12274_),
    .A2(_12277_),
    .B1(_00307_),
    .B2(_12279_),
    .C1(_12280_),
    .Y(_00042_));
 sky130_vsdinv _16382_ (.A(mem_la_wdata[0]),
    .Y(_12281_));
 sky130_fd_sc_hd__nor2_2 _16383_ (.A(_12281_),
    .B(pcpi_rs1[0]),
    .Y(_12282_));
 sky130_fd_sc_hd__or2_2 _16384_ (.A(_00048_),
    .B(_12282_),
    .X(_02591_));
 sky130_fd_sc_hd__nor2_2 _16385_ (.A(_11339_),
    .B(_11829_),
    .Y(_12283_));
 sky130_fd_sc_hd__a21oi_2 _16386_ (.A1(_11339_),
    .A2(_11829_),
    .B1(_12283_),
    .Y(_12284_));
 sky130_fd_sc_hd__nor2_2 _16387_ (.A(_11340_),
    .B(_11831_),
    .Y(_12285_));
 sky130_fd_sc_hd__a21oi_2 _16388_ (.A1(_11340_),
    .A2(_11831_),
    .B1(_12285_),
    .Y(_12286_));
 sky130_fd_sc_hd__nor2_2 _16389_ (.A(pcpi_rs2[22]),
    .B(_11830_),
    .Y(_12287_));
 sky130_fd_sc_hd__a21oi_2 _16390_ (.A1(pcpi_rs2[22]),
    .A2(_11830_),
    .B1(_12287_),
    .Y(_12288_));
 sky130_fd_sc_hd__nor2_2 _16391_ (.A(pcpi_rs2[20]),
    .B(_11832_),
    .Y(_12289_));
 sky130_fd_sc_hd__a21oi_2 _16392_ (.A1(pcpi_rs2[20]),
    .A2(_11832_),
    .B1(_12289_),
    .Y(_12290_));
 sky130_fd_sc_hd__or4_2 _16393_ (.A(_12284_),
    .B(_12286_),
    .C(_12288_),
    .D(_12290_),
    .X(_12291_));
 sky130_fd_sc_hd__nor2_2 _16394_ (.A(pcpi_rs2[16]),
    .B(_11839_),
    .Y(_12292_));
 sky130_fd_sc_hd__a21oi_2 _16395_ (.A1(pcpi_rs2[16]),
    .A2(_11839_),
    .B1(_12292_),
    .Y(_12293_));
 sky130_fd_sc_hd__nor2_2 _16396_ (.A(pcpi_rs2[18]),
    .B(_11836_),
    .Y(_12294_));
 sky130_fd_sc_hd__a21oi_2 _16397_ (.A1(pcpi_rs2[18]),
    .A2(_11836_),
    .B1(_12294_),
    .Y(_12295_));
 sky130_fd_sc_hd__nor2_2 _16398_ (.A(_11344_),
    .B(_11838_),
    .Y(_12296_));
 sky130_fd_sc_hd__a21oi_2 _16399_ (.A1(_11344_),
    .A2(_11838_),
    .B1(_12296_),
    .Y(_12297_));
 sky130_fd_sc_hd__nor2_2 _16400_ (.A(_11342_),
    .B(_11834_),
    .Y(_12298_));
 sky130_fd_sc_hd__a21oi_2 _16401_ (.A1(_11342_),
    .A2(_11834_),
    .B1(_12298_),
    .Y(_12299_));
 sky130_fd_sc_hd__or4_2 _16402_ (.A(_12293_),
    .B(_12295_),
    .C(_12297_),
    .D(_12299_),
    .X(_12300_));
 sky130_fd_sc_hd__nor2_2 _16403_ (.A(pcpi_rs2[29]),
    .B(pcpi_rs1[29]),
    .Y(_12301_));
 sky130_fd_sc_hd__a21oi_2 _16404_ (.A1(_11334_),
    .A2(pcpi_rs1[29]),
    .B1(_12301_),
    .Y(_12302_));
 sky130_fd_sc_hd__nor2_2 _16405_ (.A(pcpi_rs2[28]),
    .B(pcpi_rs1[28]),
    .Y(_12303_));
 sky130_fd_sc_hd__a21oi_2 _16406_ (.A1(pcpi_rs2[28]),
    .A2(pcpi_rs1[28]),
    .B1(_12303_),
    .Y(_12304_));
 sky130_fd_sc_hd__nor2_2 _16407_ (.A(pcpi_rs1[31]),
    .B(pcpi_rs2[31]),
    .Y(_12305_));
 sky130_fd_sc_hd__a21oi_2 _16408_ (.A1(pcpi_rs1[31]),
    .A2(pcpi_rs2[31]),
    .B1(_12305_),
    .Y(_12306_));
 sky130_fd_sc_hd__nor2_2 _16409_ (.A(pcpi_rs2[30]),
    .B(pcpi_rs1[30]),
    .Y(_12307_));
 sky130_fd_sc_hd__a21oi_2 _16410_ (.A1(pcpi_rs2[30]),
    .A2(pcpi_rs1[30]),
    .B1(_12307_),
    .Y(_12308_));
 sky130_fd_sc_hd__or2_2 _16411_ (.A(_12306_),
    .B(_12308_),
    .X(_12309_));
 sky130_fd_sc_hd__nor2_2 _16412_ (.A(pcpi_rs2[27]),
    .B(pcpi_rs1[27]),
    .Y(_12310_));
 sky130_fd_sc_hd__a21oi_2 _16413_ (.A1(_11335_),
    .A2(_11819_),
    .B1(_12310_),
    .Y(_12311_));
 sky130_fd_sc_hd__nor2_2 _16414_ (.A(pcpi_rs2[26]),
    .B(pcpi_rs1[26]),
    .Y(_12312_));
 sky130_fd_sc_hd__a21oi_2 _16415_ (.A1(pcpi_rs2[26]),
    .A2(_11821_),
    .B1(_12312_),
    .Y(_12313_));
 sky130_fd_sc_hd__nor2_2 _16416_ (.A(pcpi_rs2[25]),
    .B(pcpi_rs1[25]),
    .Y(_12314_));
 sky130_fd_sc_hd__a21oi_2 _16417_ (.A1(_11337_),
    .A2(_11824_),
    .B1(_12314_),
    .Y(_12315_));
 sky130_fd_sc_hd__nor2_2 _16418_ (.A(pcpi_rs2[24]),
    .B(_11828_),
    .Y(_12316_));
 sky130_fd_sc_hd__a21oi_2 _16419_ (.A1(pcpi_rs2[24]),
    .A2(_11828_),
    .B1(_12316_),
    .Y(_12317_));
 sky130_fd_sc_hd__or4_2 _16420_ (.A(_12311_),
    .B(_12313_),
    .C(_12315_),
    .D(_12317_),
    .X(_12318_));
 sky130_fd_sc_hd__or4_2 _16421_ (.A(_12302_),
    .B(_12304_),
    .C(_12309_),
    .D(_12318_),
    .X(_12319_));
 sky130_fd_sc_hd__nor2_2 _16422_ (.A(mem_la_wdata[5]),
    .B(pcpi_rs1[5]),
    .Y(_12320_));
 sky130_fd_sc_hd__a21oi_2 _16423_ (.A1(_11359_),
    .A2(_11857_),
    .B1(_12320_),
    .Y(_12321_));
 sky130_fd_sc_hd__nor2_2 _16424_ (.A(mem_la_wdata[7]),
    .B(_11853_),
    .Y(_12322_));
 sky130_fd_sc_hd__a21oi_2 _16425_ (.A1(_11356_),
    .A2(_11853_),
    .B1(_12322_),
    .Y(_12323_));
 sky130_fd_sc_hd__nor2_2 _16426_ (.A(_11363_),
    .B(_11862_),
    .Y(_12324_));
 sky130_fd_sc_hd__a21oi_2 _16427_ (.A1(_11363_),
    .A2(_11862_),
    .B1(_12324_),
    .Y(_12325_));
 sky130_fd_sc_hd__nor2_2 _16428_ (.A(mem_la_wdata[3]),
    .B(pcpi_rs1[3]),
    .Y(_12326_));
 sky130_fd_sc_hd__a21oi_2 _16429_ (.A1(_11361_),
    .A2(_11859_),
    .B1(_12326_),
    .Y(_12327_));
 sky130_fd_sc_hd__or4_2 _16430_ (.A(_12321_),
    .B(_12323_),
    .C(_12325_),
    .D(_12327_),
    .X(_12328_));
 sky130_fd_sc_hd__nor2_2 _16431_ (.A(mem_la_wdata[4]),
    .B(pcpi_rs1[4]),
    .Y(_12329_));
 sky130_fd_sc_hd__a21oi_2 _16432_ (.A1(_11360_),
    .A2(_11858_),
    .B1(_12329_),
    .Y(_12330_));
 sky130_fd_sc_hd__nor2_2 _16433_ (.A(mem_la_wdata[6]),
    .B(_11855_),
    .Y(_12331_));
 sky130_fd_sc_hd__a21oi_2 _16434_ (.A1(_11358_),
    .A2(_11856_),
    .B1(_12331_),
    .Y(_12332_));
 sky130_fd_sc_hd__nor2_2 _16435_ (.A(mem_la_wdata[2]),
    .B(pcpi_rs1[2]),
    .Y(_12333_));
 sky130_fd_sc_hd__a21oi_2 _16436_ (.A1(mem_la_wdata[2]),
    .A2(_11860_),
    .B1(_12333_),
    .Y(_12334_));
 sky130_fd_sc_hd__or4_2 _16437_ (.A(_02591_),
    .B(_12330_),
    .C(_12332_),
    .D(_12334_),
    .X(_12335_));
 sky130_fd_sc_hd__nor2_2 _16438_ (.A(pcpi_rs2[15]),
    .B(_11840_),
    .Y(_12336_));
 sky130_fd_sc_hd__a21oi_2 _16439_ (.A1(_11345_),
    .A2(_11840_),
    .B1(_12336_),
    .Y(_12337_));
 sky130_fd_sc_hd__nor2_2 _16440_ (.A(_11350_),
    .B(_11845_),
    .Y(_12338_));
 sky130_fd_sc_hd__a21oi_2 _16441_ (.A1(_11350_),
    .A2(_11845_),
    .B1(_12338_),
    .Y(_12339_));
 sky130_fd_sc_hd__nor2_2 _16442_ (.A(pcpi_rs2[13]),
    .B(_11843_),
    .Y(_12340_));
 sky130_fd_sc_hd__a21oi_2 _16443_ (.A1(_11348_),
    .A2(_11843_),
    .B1(_12340_),
    .Y(_12341_));
 sky130_fd_sc_hd__nor2_2 _16444_ (.A(_11346_),
    .B(_11841_),
    .Y(_12342_));
 sky130_fd_sc_hd__a21oi_2 _16445_ (.A1(_11346_),
    .A2(_11841_),
    .B1(_12342_),
    .Y(_12343_));
 sky130_fd_sc_hd__or4_2 _16446_ (.A(_12337_),
    .B(_12339_),
    .C(_12341_),
    .D(_12343_),
    .X(_12344_));
 sky130_fd_sc_hd__nor2_2 _16447_ (.A(pcpi_rs2[11]),
    .B(_11846_),
    .Y(_12345_));
 sky130_fd_sc_hd__a21oi_2 _16448_ (.A1(_11351_),
    .A2(_11846_),
    .B1(_12345_),
    .Y(_12346_));
 sky130_fd_sc_hd__nor2_2 _16449_ (.A(_11354_),
    .B(_11850_),
    .Y(_12347_));
 sky130_fd_sc_hd__a21oi_2 _16450_ (.A1(_11354_),
    .A2(_11850_),
    .B1(_12347_),
    .Y(_12348_));
 sky130_fd_sc_hd__nor2_2 _16451_ (.A(pcpi_rs2[9]),
    .B(_11849_),
    .Y(_12349_));
 sky130_fd_sc_hd__a21oi_2 _16452_ (.A1(_11353_),
    .A2(_11849_),
    .B1(_12349_),
    .Y(_12350_));
 sky130_fd_sc_hd__nor2_2 _16453_ (.A(_11352_),
    .B(_11847_),
    .Y(_12351_));
 sky130_fd_sc_hd__a21oi_2 _16454_ (.A1(_11352_),
    .A2(_11847_),
    .B1(_12351_),
    .Y(_12352_));
 sky130_fd_sc_hd__or4_2 _16455_ (.A(_12346_),
    .B(_12348_),
    .C(_12350_),
    .D(_12352_),
    .X(_12353_));
 sky130_fd_sc_hd__or4_2 _16456_ (.A(_12328_),
    .B(_12335_),
    .C(_12344_),
    .D(_12353_),
    .X(_12354_));
 sky130_fd_sc_hd__or4_2 _16457_ (.A(_12291_),
    .B(_12300_),
    .C(_12319_),
    .D(_12354_),
    .X(_12355_));
 sky130_fd_sc_hd__inv_2 _16458_ (.A(_12355_),
    .Y(_00000_));
 sky130_fd_sc_hd__or2_2 _16459_ (.A(_10581_),
    .B(_10582_),
    .X(\pcpi_mul.instr_any_mulh ));
 sky130_fd_sc_hd__or3_2 _16460_ (.A(instr_slt),
    .B(instr_slti),
    .C(instr_blt),
    .X(_00006_));
 sky130_fd_sc_hd__or3_2 _16461_ (.A(instr_sltu),
    .B(instr_sltiu),
    .C(instr_bltu),
    .X(_00007_));
 sky130_fd_sc_hd__or2_2 _16462_ (.A(mem_xfer),
    .B(_10478_),
    .X(_00299_));
 sky130_vsdinv _16463_ (.A(instr_sh),
    .Y(_12356_));
 sky130_fd_sc_hd__nor2_2 _16464_ (.A(instr_lhu),
    .B(instr_lh),
    .Y(_12357_));
 sky130_fd_sc_hd__o32a_2 _16465_ (.A1(_12356_),
    .A2(_11807_),
    .A3(_10809_),
    .B1(_10812_),
    .B2(_12357_),
    .X(_12358_));
 sky130_fd_sc_hd__buf_1 _16466_ (.A(_12207_),
    .X(_12359_));
 sky130_fd_sc_hd__buf_1 _16467_ (.A(_12359_),
    .X(_12360_));
 sky130_fd_sc_hd__nor2_2 _16468_ (.A(_00319_),
    .B(_00317_),
    .Y(_12361_));
 sky130_fd_sc_hd__o21a_2 _16469_ (.A1(_10651_),
    .A2(_10671_),
    .B1(_10443_),
    .X(_12362_));
 sky130_fd_sc_hd__o221a_2 _16470_ (.A1(_00297_),
    .A2(_12258_),
    .B1(_00296_),
    .B2(_12361_),
    .C1(_12362_),
    .X(_12363_));
 sky130_fd_sc_hd__o22ai_2 _16471_ (.A1(_00296_),
    .A2(_12358_),
    .B1(_12360_),
    .B2(_12363_),
    .Y(_00047_));
 sky130_fd_sc_hd__buf_1 _16472_ (.A(_10604_),
    .X(_12364_));
 sky130_fd_sc_hd__nor2_2 _16473_ (.A(_12364_),
    .B(_10671_),
    .Y(_00336_));
 sky130_fd_sc_hd__nor2_2 _16474_ (.A(_12947_),
    .B(_12260_),
    .Y(_00338_));
 sky130_vsdinv _16475_ (.A(alu_eq),
    .Y(_00340_));
 sky130_fd_sc_hd__or3_2 _16476_ (.A(instr_bne),
    .B(is_slti_blt_slt),
    .C(is_sltiu_bltu_sltu),
    .X(_12365_));
 sky130_fd_sc_hd__nor3_2 _16477_ (.A(instr_bgeu),
    .B(instr_bge),
    .C(_12365_),
    .Y(_00341_));
 sky130_fd_sc_hd__mux2_2 _16478_ (.A0(instr_bgeu),
    .A1(is_sltiu_bltu_sltu),
    .S(alu_ltu),
    .X(_12366_));
 sky130_fd_sc_hd__a21oi_2 _16479_ (.A1(is_slti_blt_slt),
    .A2(alu_lts),
    .B1(_12366_),
    .Y(_12367_));
 sky130_fd_sc_hd__o221a_2 _16480_ (.A1(_10798_),
    .A2(alu_eq),
    .B1(_10794_),
    .B2(alu_lts),
    .C1(_12367_),
    .X(_00342_));
 sky130_vsdinv _16481_ (.A(_00343_),
    .Y(_12368_));
 sky130_fd_sc_hd__or2_2 _16482_ (.A(_12368_),
    .B(_00337_),
    .X(_00344_));
 sky130_fd_sc_hd__o22ai_2 _16483_ (.A1(_00339_),
    .A2(_00297_),
    .B1(_12274_),
    .B2(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__o21a_2 _16484_ (.A1(decoder_trigger),
    .A2(do_waitirq),
    .B1(_10648_),
    .X(_00349_));
 sky130_fd_sc_hd__and2_2 _16485_ (.A(_02410_),
    .B(_00349_),
    .X(_00351_));
 sky130_fd_sc_hd__and3_2 _16486_ (.A(_11030_),
    .B(_12182_),
    .C(_10609_),
    .X(_00354_));
 sky130_fd_sc_hd__buf_1 _16487_ (.A(_11080_),
    .X(_12369_));
 sky130_fd_sc_hd__o211a_2 _16488_ (.A1(_12274_),
    .A2(_12257_),
    .B1(_12369_),
    .C1(_12182_),
    .X(_00355_));
 sky130_vsdinv _16489_ (.A(\cpuregs[0][1] ),
    .Y(_00371_));
 sky130_vsdinv _16490_ (.A(\cpuregs[1][1] ),
    .Y(_00372_));
 sky130_vsdinv _16491_ (.A(\cpuregs[2][1] ),
    .Y(_00373_));
 sky130_vsdinv _16492_ (.A(\cpuregs[3][1] ),
    .Y(_00374_));
 sky130_vsdinv _16493_ (.A(\cpuregs[4][1] ),
    .Y(_00376_));
 sky130_vsdinv _16494_ (.A(\cpuregs[5][1] ),
    .Y(_00377_));
 sky130_vsdinv _16495_ (.A(\cpuregs[6][1] ),
    .Y(_00378_));
 sky130_vsdinv _16496_ (.A(\cpuregs[7][1] ),
    .Y(_00379_));
 sky130_vsdinv _16497_ (.A(\cpuregs[8][1] ),
    .Y(_00381_));
 sky130_vsdinv _16498_ (.A(\cpuregs[9][1] ),
    .Y(_00382_));
 sky130_vsdinv _16499_ (.A(\cpuregs[10][1] ),
    .Y(_00383_));
 sky130_vsdinv _16500_ (.A(\cpuregs[11][1] ),
    .Y(_00384_));
 sky130_vsdinv _16501_ (.A(\cpuregs[12][1] ),
    .Y(_00386_));
 sky130_vsdinv _16502_ (.A(\cpuregs[13][1] ),
    .Y(_00387_));
 sky130_vsdinv _16503_ (.A(\cpuregs[14][1] ),
    .Y(_00388_));
 sky130_vsdinv _16504_ (.A(\cpuregs[15][1] ),
    .Y(_00389_));
 sky130_vsdinv _16505_ (.A(\cpuregs[16][1] ),
    .Y(_00392_));
 sky130_vsdinv _16506_ (.A(\cpuregs[17][1] ),
    .Y(_00393_));
 sky130_vsdinv _16507_ (.A(\cpuregs[18][1] ),
    .Y(_00394_));
 sky130_vsdinv _16508_ (.A(\cpuregs[19][1] ),
    .Y(_00395_));
 sky130_vsdinv _16509_ (.A(\cpuregs[0][2] ),
    .Y(_00398_));
 sky130_vsdinv _16510_ (.A(\cpuregs[1][2] ),
    .Y(_00399_));
 sky130_vsdinv _16511_ (.A(\cpuregs[2][2] ),
    .Y(_00400_));
 sky130_vsdinv _16512_ (.A(\cpuregs[3][2] ),
    .Y(_00401_));
 sky130_vsdinv _16513_ (.A(\cpuregs[4][2] ),
    .Y(_00403_));
 sky130_vsdinv _16514_ (.A(\cpuregs[5][2] ),
    .Y(_00404_));
 sky130_vsdinv _16515_ (.A(\cpuregs[6][2] ),
    .Y(_00405_));
 sky130_vsdinv _16516_ (.A(\cpuregs[7][2] ),
    .Y(_00406_));
 sky130_vsdinv _16517_ (.A(\cpuregs[8][2] ),
    .Y(_00408_));
 sky130_vsdinv _16518_ (.A(\cpuregs[9][2] ),
    .Y(_00409_));
 sky130_vsdinv _16519_ (.A(\cpuregs[10][2] ),
    .Y(_00410_));
 sky130_vsdinv _16520_ (.A(\cpuregs[11][2] ),
    .Y(_00411_));
 sky130_vsdinv _16521_ (.A(\cpuregs[12][2] ),
    .Y(_00413_));
 sky130_vsdinv _16522_ (.A(\cpuregs[13][2] ),
    .Y(_00414_));
 sky130_vsdinv _16523_ (.A(\cpuregs[14][2] ),
    .Y(_00415_));
 sky130_vsdinv _16524_ (.A(\cpuregs[15][2] ),
    .Y(_00416_));
 sky130_vsdinv _16525_ (.A(\cpuregs[16][2] ),
    .Y(_00419_));
 sky130_vsdinv _16526_ (.A(\cpuregs[17][2] ),
    .Y(_00420_));
 sky130_vsdinv _16527_ (.A(\cpuregs[18][2] ),
    .Y(_00421_));
 sky130_vsdinv _16528_ (.A(\cpuregs[19][2] ),
    .Y(_00422_));
 sky130_vsdinv _16529_ (.A(\cpuregs[0][3] ),
    .Y(_00425_));
 sky130_vsdinv _16530_ (.A(\cpuregs[1][3] ),
    .Y(_00426_));
 sky130_vsdinv _16531_ (.A(\cpuregs[2][3] ),
    .Y(_00427_));
 sky130_vsdinv _16532_ (.A(\cpuregs[3][3] ),
    .Y(_00428_));
 sky130_vsdinv _16533_ (.A(\cpuregs[4][3] ),
    .Y(_00430_));
 sky130_vsdinv _16534_ (.A(\cpuregs[5][3] ),
    .Y(_00431_));
 sky130_vsdinv _16535_ (.A(\cpuregs[6][3] ),
    .Y(_00432_));
 sky130_vsdinv _16536_ (.A(\cpuregs[7][3] ),
    .Y(_00433_));
 sky130_vsdinv _16537_ (.A(\cpuregs[8][3] ),
    .Y(_00435_));
 sky130_vsdinv _16538_ (.A(\cpuregs[9][3] ),
    .Y(_00436_));
 sky130_vsdinv _16539_ (.A(\cpuregs[10][3] ),
    .Y(_00437_));
 sky130_vsdinv _16540_ (.A(\cpuregs[11][3] ),
    .Y(_00438_));
 sky130_vsdinv _16541_ (.A(\cpuregs[12][3] ),
    .Y(_00440_));
 sky130_vsdinv _16542_ (.A(\cpuregs[13][3] ),
    .Y(_00441_));
 sky130_vsdinv _16543_ (.A(\cpuregs[14][3] ),
    .Y(_00442_));
 sky130_vsdinv _16544_ (.A(\cpuregs[15][3] ),
    .Y(_00443_));
 sky130_vsdinv _16545_ (.A(\cpuregs[16][3] ),
    .Y(_00446_));
 sky130_vsdinv _16546_ (.A(\cpuregs[17][3] ),
    .Y(_00447_));
 sky130_vsdinv _16547_ (.A(\cpuregs[18][3] ),
    .Y(_00448_));
 sky130_vsdinv _16548_ (.A(\cpuregs[19][3] ),
    .Y(_00449_));
 sky130_vsdinv _16549_ (.A(\cpuregs[0][4] ),
    .Y(_00452_));
 sky130_vsdinv _16550_ (.A(\cpuregs[1][4] ),
    .Y(_00453_));
 sky130_vsdinv _16551_ (.A(\cpuregs[2][4] ),
    .Y(_00454_));
 sky130_vsdinv _16552_ (.A(\cpuregs[3][4] ),
    .Y(_00455_));
 sky130_vsdinv _16553_ (.A(\cpuregs[4][4] ),
    .Y(_00457_));
 sky130_vsdinv _16554_ (.A(\cpuregs[5][4] ),
    .Y(_00458_));
 sky130_vsdinv _16555_ (.A(\cpuregs[6][4] ),
    .Y(_00459_));
 sky130_vsdinv _16556_ (.A(\cpuregs[7][4] ),
    .Y(_00460_));
 sky130_vsdinv _16557_ (.A(\cpuregs[8][4] ),
    .Y(_00462_));
 sky130_vsdinv _16558_ (.A(\cpuregs[9][4] ),
    .Y(_00463_));
 sky130_vsdinv _16559_ (.A(\cpuregs[10][4] ),
    .Y(_00464_));
 sky130_vsdinv _16560_ (.A(\cpuregs[11][4] ),
    .Y(_00465_));
 sky130_vsdinv _16561_ (.A(\cpuregs[12][4] ),
    .Y(_00467_));
 sky130_vsdinv _16562_ (.A(\cpuregs[13][4] ),
    .Y(_00468_));
 sky130_vsdinv _16563_ (.A(\cpuregs[14][4] ),
    .Y(_00469_));
 sky130_vsdinv _16564_ (.A(\cpuregs[15][4] ),
    .Y(_00470_));
 sky130_vsdinv _16565_ (.A(\cpuregs[16][4] ),
    .Y(_00473_));
 sky130_vsdinv _16566_ (.A(\cpuregs[17][4] ),
    .Y(_00474_));
 sky130_vsdinv _16567_ (.A(\cpuregs[18][4] ),
    .Y(_00475_));
 sky130_vsdinv _16568_ (.A(\cpuregs[19][4] ),
    .Y(_00476_));
 sky130_vsdinv _16569_ (.A(\cpuregs[0][5] ),
    .Y(_00479_));
 sky130_vsdinv _16570_ (.A(\cpuregs[1][5] ),
    .Y(_00480_));
 sky130_vsdinv _16571_ (.A(\cpuregs[2][5] ),
    .Y(_00481_));
 sky130_vsdinv _16572_ (.A(\cpuregs[3][5] ),
    .Y(_00482_));
 sky130_vsdinv _16573_ (.A(\cpuregs[4][5] ),
    .Y(_00484_));
 sky130_vsdinv _16574_ (.A(\cpuregs[5][5] ),
    .Y(_00485_));
 sky130_vsdinv _16575_ (.A(\cpuregs[6][5] ),
    .Y(_00486_));
 sky130_vsdinv _16576_ (.A(\cpuregs[7][5] ),
    .Y(_00487_));
 sky130_vsdinv _16577_ (.A(\cpuregs[8][5] ),
    .Y(_00489_));
 sky130_vsdinv _16578_ (.A(\cpuregs[9][5] ),
    .Y(_00490_));
 sky130_vsdinv _16579_ (.A(\cpuregs[10][5] ),
    .Y(_00491_));
 sky130_vsdinv _16580_ (.A(\cpuregs[11][5] ),
    .Y(_00492_));
 sky130_vsdinv _16581_ (.A(\cpuregs[12][5] ),
    .Y(_00494_));
 sky130_vsdinv _16582_ (.A(\cpuregs[13][5] ),
    .Y(_00495_));
 sky130_vsdinv _16583_ (.A(\cpuregs[14][5] ),
    .Y(_00496_));
 sky130_vsdinv _16584_ (.A(\cpuregs[15][5] ),
    .Y(_00497_));
 sky130_vsdinv _16585_ (.A(\cpuregs[16][5] ),
    .Y(_00500_));
 sky130_vsdinv _16586_ (.A(\cpuregs[17][5] ),
    .Y(_00501_));
 sky130_vsdinv _16587_ (.A(\cpuregs[18][5] ),
    .Y(_00502_));
 sky130_vsdinv _16588_ (.A(\cpuregs[19][5] ),
    .Y(_00503_));
 sky130_vsdinv _16589_ (.A(\cpuregs[0][6] ),
    .Y(_00506_));
 sky130_vsdinv _16590_ (.A(\cpuregs[1][6] ),
    .Y(_00507_));
 sky130_vsdinv _16591_ (.A(\cpuregs[2][6] ),
    .Y(_00508_));
 sky130_vsdinv _16592_ (.A(\cpuregs[3][6] ),
    .Y(_00509_));
 sky130_vsdinv _16593_ (.A(\cpuregs[4][6] ),
    .Y(_00511_));
 sky130_vsdinv _16594_ (.A(\cpuregs[5][6] ),
    .Y(_00512_));
 sky130_vsdinv _16595_ (.A(\cpuregs[6][6] ),
    .Y(_00513_));
 sky130_vsdinv _16596_ (.A(\cpuregs[7][6] ),
    .Y(_00514_));
 sky130_vsdinv _16597_ (.A(\cpuregs[8][6] ),
    .Y(_00516_));
 sky130_vsdinv _16598_ (.A(\cpuregs[9][6] ),
    .Y(_00517_));
 sky130_vsdinv _16599_ (.A(\cpuregs[10][6] ),
    .Y(_00518_));
 sky130_vsdinv _16600_ (.A(\cpuregs[11][6] ),
    .Y(_00519_));
 sky130_vsdinv _16601_ (.A(\cpuregs[12][6] ),
    .Y(_00521_));
 sky130_vsdinv _16602_ (.A(\cpuregs[13][6] ),
    .Y(_00522_));
 sky130_vsdinv _16603_ (.A(\cpuregs[14][6] ),
    .Y(_00523_));
 sky130_vsdinv _16604_ (.A(\cpuregs[15][6] ),
    .Y(_00524_));
 sky130_vsdinv _16605_ (.A(\cpuregs[16][6] ),
    .Y(_00527_));
 sky130_vsdinv _16606_ (.A(\cpuregs[17][6] ),
    .Y(_00528_));
 sky130_vsdinv _16607_ (.A(\cpuregs[18][6] ),
    .Y(_00529_));
 sky130_vsdinv _16608_ (.A(\cpuregs[19][6] ),
    .Y(_00530_));
 sky130_vsdinv _16609_ (.A(\cpuregs[0][7] ),
    .Y(_00533_));
 sky130_vsdinv _16610_ (.A(\cpuregs[1][7] ),
    .Y(_00534_));
 sky130_vsdinv _16611_ (.A(\cpuregs[2][7] ),
    .Y(_00535_));
 sky130_vsdinv _16612_ (.A(\cpuregs[3][7] ),
    .Y(_00536_));
 sky130_vsdinv _16613_ (.A(\cpuregs[4][7] ),
    .Y(_00538_));
 sky130_vsdinv _16614_ (.A(\cpuregs[5][7] ),
    .Y(_00539_));
 sky130_vsdinv _16615_ (.A(\cpuregs[6][7] ),
    .Y(_00540_));
 sky130_vsdinv _16616_ (.A(\cpuregs[7][7] ),
    .Y(_00541_));
 sky130_vsdinv _16617_ (.A(\cpuregs[8][7] ),
    .Y(_00543_));
 sky130_vsdinv _16618_ (.A(\cpuregs[9][7] ),
    .Y(_00544_));
 sky130_vsdinv _16619_ (.A(\cpuregs[10][7] ),
    .Y(_00545_));
 sky130_vsdinv _16620_ (.A(\cpuregs[11][7] ),
    .Y(_00546_));
 sky130_vsdinv _16621_ (.A(\cpuregs[12][7] ),
    .Y(_00548_));
 sky130_vsdinv _16622_ (.A(\cpuregs[13][7] ),
    .Y(_00549_));
 sky130_vsdinv _16623_ (.A(\cpuregs[14][7] ),
    .Y(_00550_));
 sky130_vsdinv _16624_ (.A(\cpuregs[15][7] ),
    .Y(_00551_));
 sky130_vsdinv _16625_ (.A(\cpuregs[16][7] ),
    .Y(_00554_));
 sky130_vsdinv _16626_ (.A(\cpuregs[17][7] ),
    .Y(_00555_));
 sky130_vsdinv _16627_ (.A(\cpuregs[18][7] ),
    .Y(_00556_));
 sky130_vsdinv _16628_ (.A(\cpuregs[19][7] ),
    .Y(_00557_));
 sky130_vsdinv _16629_ (.A(\cpuregs[0][8] ),
    .Y(_00560_));
 sky130_vsdinv _16630_ (.A(\cpuregs[1][8] ),
    .Y(_00561_));
 sky130_vsdinv _16631_ (.A(\cpuregs[2][8] ),
    .Y(_00562_));
 sky130_vsdinv _16632_ (.A(\cpuregs[3][8] ),
    .Y(_00563_));
 sky130_vsdinv _16633_ (.A(\cpuregs[4][8] ),
    .Y(_00565_));
 sky130_vsdinv _16634_ (.A(\cpuregs[5][8] ),
    .Y(_00566_));
 sky130_vsdinv _16635_ (.A(\cpuregs[6][8] ),
    .Y(_00567_));
 sky130_vsdinv _16636_ (.A(\cpuregs[7][8] ),
    .Y(_00568_));
 sky130_vsdinv _16637_ (.A(\cpuregs[8][8] ),
    .Y(_00570_));
 sky130_vsdinv _16638_ (.A(\cpuregs[9][8] ),
    .Y(_00571_));
 sky130_vsdinv _16639_ (.A(\cpuregs[10][8] ),
    .Y(_00572_));
 sky130_vsdinv _16640_ (.A(\cpuregs[11][8] ),
    .Y(_00573_));
 sky130_vsdinv _16641_ (.A(\cpuregs[12][8] ),
    .Y(_00575_));
 sky130_vsdinv _16642_ (.A(\cpuregs[13][8] ),
    .Y(_00576_));
 sky130_vsdinv _16643_ (.A(\cpuregs[14][8] ),
    .Y(_00577_));
 sky130_vsdinv _16644_ (.A(\cpuregs[15][8] ),
    .Y(_00578_));
 sky130_vsdinv _16645_ (.A(\cpuregs[16][8] ),
    .Y(_00581_));
 sky130_vsdinv _16646_ (.A(\cpuregs[17][8] ),
    .Y(_00582_));
 sky130_vsdinv _16647_ (.A(\cpuregs[18][8] ),
    .Y(_00583_));
 sky130_vsdinv _16648_ (.A(\cpuregs[19][8] ),
    .Y(_00584_));
 sky130_vsdinv _16649_ (.A(\cpuregs[0][9] ),
    .Y(_00587_));
 sky130_vsdinv _16650_ (.A(\cpuregs[1][9] ),
    .Y(_00588_));
 sky130_vsdinv _16651_ (.A(\cpuregs[2][9] ),
    .Y(_00589_));
 sky130_vsdinv _16652_ (.A(\cpuregs[3][9] ),
    .Y(_00590_));
 sky130_vsdinv _16653_ (.A(\cpuregs[4][9] ),
    .Y(_00592_));
 sky130_vsdinv _16654_ (.A(\cpuregs[5][9] ),
    .Y(_00593_));
 sky130_vsdinv _16655_ (.A(\cpuregs[6][9] ),
    .Y(_00594_));
 sky130_vsdinv _16656_ (.A(\cpuregs[7][9] ),
    .Y(_00595_));
 sky130_vsdinv _16657_ (.A(\cpuregs[8][9] ),
    .Y(_00597_));
 sky130_vsdinv _16658_ (.A(\cpuregs[9][9] ),
    .Y(_00598_));
 sky130_vsdinv _16659_ (.A(\cpuregs[10][9] ),
    .Y(_00599_));
 sky130_vsdinv _16660_ (.A(\cpuregs[11][9] ),
    .Y(_00600_));
 sky130_vsdinv _16661_ (.A(\cpuregs[12][9] ),
    .Y(_00602_));
 sky130_vsdinv _16662_ (.A(\cpuregs[13][9] ),
    .Y(_00603_));
 sky130_vsdinv _16663_ (.A(\cpuregs[14][9] ),
    .Y(_00604_));
 sky130_vsdinv _16664_ (.A(\cpuregs[15][9] ),
    .Y(_00605_));
 sky130_vsdinv _16665_ (.A(\cpuregs[16][9] ),
    .Y(_00608_));
 sky130_vsdinv _16666_ (.A(\cpuregs[17][9] ),
    .Y(_00609_));
 sky130_vsdinv _16667_ (.A(\cpuregs[18][9] ),
    .Y(_00610_));
 sky130_vsdinv _16668_ (.A(\cpuregs[19][9] ),
    .Y(_00611_));
 sky130_vsdinv _16669_ (.A(\cpuregs[0][10] ),
    .Y(_00614_));
 sky130_vsdinv _16670_ (.A(\cpuregs[1][10] ),
    .Y(_00615_));
 sky130_vsdinv _16671_ (.A(\cpuregs[2][10] ),
    .Y(_00616_));
 sky130_vsdinv _16672_ (.A(\cpuregs[3][10] ),
    .Y(_00617_));
 sky130_vsdinv _16673_ (.A(\cpuregs[4][10] ),
    .Y(_00619_));
 sky130_vsdinv _16674_ (.A(\cpuregs[5][10] ),
    .Y(_00620_));
 sky130_vsdinv _16675_ (.A(\cpuregs[6][10] ),
    .Y(_00621_));
 sky130_vsdinv _16676_ (.A(\cpuregs[7][10] ),
    .Y(_00622_));
 sky130_vsdinv _16677_ (.A(\cpuregs[8][10] ),
    .Y(_00624_));
 sky130_vsdinv _16678_ (.A(\cpuregs[9][10] ),
    .Y(_00625_));
 sky130_vsdinv _16679_ (.A(\cpuregs[10][10] ),
    .Y(_00626_));
 sky130_vsdinv _16680_ (.A(\cpuregs[11][10] ),
    .Y(_00627_));
 sky130_vsdinv _16681_ (.A(\cpuregs[12][10] ),
    .Y(_00629_));
 sky130_vsdinv _16682_ (.A(\cpuregs[13][10] ),
    .Y(_00630_));
 sky130_vsdinv _16683_ (.A(\cpuregs[14][10] ),
    .Y(_00631_));
 sky130_vsdinv _16684_ (.A(\cpuregs[15][10] ),
    .Y(_00632_));
 sky130_vsdinv _16685_ (.A(\cpuregs[16][10] ),
    .Y(_00635_));
 sky130_vsdinv _16686_ (.A(\cpuregs[17][10] ),
    .Y(_00636_));
 sky130_vsdinv _16687_ (.A(\cpuregs[18][10] ),
    .Y(_00637_));
 sky130_vsdinv _16688_ (.A(\cpuregs[19][10] ),
    .Y(_00638_));
 sky130_vsdinv _16689_ (.A(\cpuregs[0][11] ),
    .Y(_00641_));
 sky130_vsdinv _16690_ (.A(\cpuregs[1][11] ),
    .Y(_00642_));
 sky130_vsdinv _16691_ (.A(\cpuregs[2][11] ),
    .Y(_00643_));
 sky130_vsdinv _16692_ (.A(\cpuregs[3][11] ),
    .Y(_00644_));
 sky130_vsdinv _16693_ (.A(\cpuregs[4][11] ),
    .Y(_00646_));
 sky130_vsdinv _16694_ (.A(\cpuregs[5][11] ),
    .Y(_00647_));
 sky130_vsdinv _16695_ (.A(\cpuregs[6][11] ),
    .Y(_00648_));
 sky130_vsdinv _16696_ (.A(\cpuregs[7][11] ),
    .Y(_00649_));
 sky130_vsdinv _16697_ (.A(\cpuregs[8][11] ),
    .Y(_00651_));
 sky130_vsdinv _16698_ (.A(\cpuregs[9][11] ),
    .Y(_00652_));
 sky130_vsdinv _16699_ (.A(\cpuregs[10][11] ),
    .Y(_00653_));
 sky130_vsdinv _16700_ (.A(\cpuregs[11][11] ),
    .Y(_00654_));
 sky130_vsdinv _16701_ (.A(\cpuregs[12][11] ),
    .Y(_00656_));
 sky130_vsdinv _16702_ (.A(\cpuregs[13][11] ),
    .Y(_00657_));
 sky130_vsdinv _16703_ (.A(\cpuregs[14][11] ),
    .Y(_00658_));
 sky130_vsdinv _16704_ (.A(\cpuregs[15][11] ),
    .Y(_00659_));
 sky130_vsdinv _16705_ (.A(\cpuregs[16][11] ),
    .Y(_00662_));
 sky130_vsdinv _16706_ (.A(\cpuregs[17][11] ),
    .Y(_00663_));
 sky130_vsdinv _16707_ (.A(\cpuregs[18][11] ),
    .Y(_00664_));
 sky130_vsdinv _16708_ (.A(\cpuregs[19][11] ),
    .Y(_00665_));
 sky130_vsdinv _16709_ (.A(\cpuregs[0][12] ),
    .Y(_00668_));
 sky130_vsdinv _16710_ (.A(\cpuregs[1][12] ),
    .Y(_00669_));
 sky130_vsdinv _16711_ (.A(\cpuregs[2][12] ),
    .Y(_00670_));
 sky130_vsdinv _16712_ (.A(\cpuregs[3][12] ),
    .Y(_00671_));
 sky130_vsdinv _16713_ (.A(\cpuregs[4][12] ),
    .Y(_00673_));
 sky130_vsdinv _16714_ (.A(\cpuregs[5][12] ),
    .Y(_00674_));
 sky130_vsdinv _16715_ (.A(\cpuregs[6][12] ),
    .Y(_00675_));
 sky130_vsdinv _16716_ (.A(\cpuregs[7][12] ),
    .Y(_00676_));
 sky130_vsdinv _16717_ (.A(\cpuregs[8][12] ),
    .Y(_00678_));
 sky130_vsdinv _16718_ (.A(\cpuregs[9][12] ),
    .Y(_00679_));
 sky130_vsdinv _16719_ (.A(\cpuregs[10][12] ),
    .Y(_00680_));
 sky130_vsdinv _16720_ (.A(\cpuregs[11][12] ),
    .Y(_00681_));
 sky130_vsdinv _16721_ (.A(\cpuregs[12][12] ),
    .Y(_00683_));
 sky130_vsdinv _16722_ (.A(\cpuregs[13][12] ),
    .Y(_00684_));
 sky130_vsdinv _16723_ (.A(\cpuregs[14][12] ),
    .Y(_00685_));
 sky130_vsdinv _16724_ (.A(\cpuregs[15][12] ),
    .Y(_00686_));
 sky130_vsdinv _16725_ (.A(\cpuregs[16][12] ),
    .Y(_00689_));
 sky130_vsdinv _16726_ (.A(\cpuregs[17][12] ),
    .Y(_00690_));
 sky130_vsdinv _16727_ (.A(\cpuregs[18][12] ),
    .Y(_00691_));
 sky130_vsdinv _16728_ (.A(\cpuregs[19][12] ),
    .Y(_00692_));
 sky130_vsdinv _16729_ (.A(\cpuregs[0][13] ),
    .Y(_00695_));
 sky130_vsdinv _16730_ (.A(\cpuregs[1][13] ),
    .Y(_00696_));
 sky130_vsdinv _16731_ (.A(\cpuregs[2][13] ),
    .Y(_00697_));
 sky130_vsdinv _16732_ (.A(\cpuregs[3][13] ),
    .Y(_00698_));
 sky130_vsdinv _16733_ (.A(\cpuregs[4][13] ),
    .Y(_00700_));
 sky130_vsdinv _16734_ (.A(\cpuregs[5][13] ),
    .Y(_00701_));
 sky130_vsdinv _16735_ (.A(\cpuregs[6][13] ),
    .Y(_00702_));
 sky130_vsdinv _16736_ (.A(\cpuregs[7][13] ),
    .Y(_00703_));
 sky130_vsdinv _16737_ (.A(\cpuregs[8][13] ),
    .Y(_00705_));
 sky130_vsdinv _16738_ (.A(\cpuregs[9][13] ),
    .Y(_00706_));
 sky130_vsdinv _16739_ (.A(\cpuregs[10][13] ),
    .Y(_00707_));
 sky130_vsdinv _16740_ (.A(\cpuregs[11][13] ),
    .Y(_00708_));
 sky130_vsdinv _16741_ (.A(\cpuregs[12][13] ),
    .Y(_00710_));
 sky130_vsdinv _16742_ (.A(\cpuregs[13][13] ),
    .Y(_00711_));
 sky130_vsdinv _16743_ (.A(\cpuregs[14][13] ),
    .Y(_00712_));
 sky130_vsdinv _16744_ (.A(\cpuregs[15][13] ),
    .Y(_00713_));
 sky130_vsdinv _16745_ (.A(\cpuregs[16][13] ),
    .Y(_00716_));
 sky130_vsdinv _16746_ (.A(\cpuregs[17][13] ),
    .Y(_00717_));
 sky130_vsdinv _16747_ (.A(\cpuregs[18][13] ),
    .Y(_00718_));
 sky130_vsdinv _16748_ (.A(\cpuregs[19][13] ),
    .Y(_00719_));
 sky130_vsdinv _16749_ (.A(\cpuregs[0][14] ),
    .Y(_00722_));
 sky130_vsdinv _16750_ (.A(\cpuregs[1][14] ),
    .Y(_00723_));
 sky130_vsdinv _16751_ (.A(\cpuregs[2][14] ),
    .Y(_00724_));
 sky130_vsdinv _16752_ (.A(\cpuregs[3][14] ),
    .Y(_00725_));
 sky130_vsdinv _16753_ (.A(\cpuregs[4][14] ),
    .Y(_00727_));
 sky130_vsdinv _16754_ (.A(\cpuregs[5][14] ),
    .Y(_00728_));
 sky130_vsdinv _16755_ (.A(\cpuregs[6][14] ),
    .Y(_00729_));
 sky130_vsdinv _16756_ (.A(\cpuregs[7][14] ),
    .Y(_00730_));
 sky130_vsdinv _16757_ (.A(\cpuregs[8][14] ),
    .Y(_00732_));
 sky130_vsdinv _16758_ (.A(\cpuregs[9][14] ),
    .Y(_00733_));
 sky130_vsdinv _16759_ (.A(\cpuregs[10][14] ),
    .Y(_00734_));
 sky130_vsdinv _16760_ (.A(\cpuregs[11][14] ),
    .Y(_00735_));
 sky130_vsdinv _16761_ (.A(\cpuregs[12][14] ),
    .Y(_00737_));
 sky130_vsdinv _16762_ (.A(\cpuregs[13][14] ),
    .Y(_00738_));
 sky130_vsdinv _16763_ (.A(\cpuregs[14][14] ),
    .Y(_00739_));
 sky130_vsdinv _16764_ (.A(\cpuregs[15][14] ),
    .Y(_00740_));
 sky130_vsdinv _16765_ (.A(\cpuregs[16][14] ),
    .Y(_00743_));
 sky130_vsdinv _16766_ (.A(\cpuregs[17][14] ),
    .Y(_00744_));
 sky130_vsdinv _16767_ (.A(\cpuregs[18][14] ),
    .Y(_00745_));
 sky130_vsdinv _16768_ (.A(\cpuregs[19][14] ),
    .Y(_00746_));
 sky130_vsdinv _16769_ (.A(\cpuregs[0][15] ),
    .Y(_00749_));
 sky130_vsdinv _16770_ (.A(\cpuregs[1][15] ),
    .Y(_00750_));
 sky130_vsdinv _16771_ (.A(\cpuregs[2][15] ),
    .Y(_00751_));
 sky130_vsdinv _16772_ (.A(\cpuregs[3][15] ),
    .Y(_00752_));
 sky130_vsdinv _16773_ (.A(\cpuregs[4][15] ),
    .Y(_00754_));
 sky130_vsdinv _16774_ (.A(\cpuregs[5][15] ),
    .Y(_00755_));
 sky130_vsdinv _16775_ (.A(\cpuregs[6][15] ),
    .Y(_00756_));
 sky130_vsdinv _16776_ (.A(\cpuregs[7][15] ),
    .Y(_00757_));
 sky130_vsdinv _16777_ (.A(\cpuregs[8][15] ),
    .Y(_00759_));
 sky130_vsdinv _16778_ (.A(\cpuregs[9][15] ),
    .Y(_00760_));
 sky130_vsdinv _16779_ (.A(\cpuregs[10][15] ),
    .Y(_00761_));
 sky130_vsdinv _16780_ (.A(\cpuregs[11][15] ),
    .Y(_00762_));
 sky130_vsdinv _16781_ (.A(\cpuregs[12][15] ),
    .Y(_00764_));
 sky130_vsdinv _16782_ (.A(\cpuregs[13][15] ),
    .Y(_00765_));
 sky130_vsdinv _16783_ (.A(\cpuregs[14][15] ),
    .Y(_00766_));
 sky130_vsdinv _16784_ (.A(\cpuregs[15][15] ),
    .Y(_00767_));
 sky130_vsdinv _16785_ (.A(\cpuregs[16][15] ),
    .Y(_00770_));
 sky130_vsdinv _16786_ (.A(\cpuregs[17][15] ),
    .Y(_00771_));
 sky130_vsdinv _16787_ (.A(\cpuregs[18][15] ),
    .Y(_00772_));
 sky130_vsdinv _16788_ (.A(\cpuregs[19][15] ),
    .Y(_00773_));
 sky130_vsdinv _16789_ (.A(\cpuregs[0][16] ),
    .Y(_00776_));
 sky130_vsdinv _16790_ (.A(\cpuregs[1][16] ),
    .Y(_00777_));
 sky130_vsdinv _16791_ (.A(\cpuregs[2][16] ),
    .Y(_00778_));
 sky130_vsdinv _16792_ (.A(\cpuregs[3][16] ),
    .Y(_00779_));
 sky130_vsdinv _16793_ (.A(\cpuregs[4][16] ),
    .Y(_00781_));
 sky130_vsdinv _16794_ (.A(\cpuregs[5][16] ),
    .Y(_00782_));
 sky130_vsdinv _16795_ (.A(\cpuregs[6][16] ),
    .Y(_00783_));
 sky130_vsdinv _16796_ (.A(\cpuregs[7][16] ),
    .Y(_00784_));
 sky130_vsdinv _16797_ (.A(\cpuregs[8][16] ),
    .Y(_00786_));
 sky130_vsdinv _16798_ (.A(\cpuregs[9][16] ),
    .Y(_00787_));
 sky130_vsdinv _16799_ (.A(\cpuregs[10][16] ),
    .Y(_00788_));
 sky130_vsdinv _16800_ (.A(\cpuregs[11][16] ),
    .Y(_00789_));
 sky130_vsdinv _16801_ (.A(\cpuregs[12][16] ),
    .Y(_00791_));
 sky130_vsdinv _16802_ (.A(\cpuregs[13][16] ),
    .Y(_00792_));
 sky130_vsdinv _16803_ (.A(\cpuregs[14][16] ),
    .Y(_00793_));
 sky130_vsdinv _16804_ (.A(\cpuregs[15][16] ),
    .Y(_00794_));
 sky130_vsdinv _16805_ (.A(\cpuregs[16][16] ),
    .Y(_00797_));
 sky130_vsdinv _16806_ (.A(\cpuregs[17][16] ),
    .Y(_00798_));
 sky130_vsdinv _16807_ (.A(\cpuregs[18][16] ),
    .Y(_00799_));
 sky130_vsdinv _16808_ (.A(\cpuregs[19][16] ),
    .Y(_00800_));
 sky130_vsdinv _16809_ (.A(\cpuregs[0][17] ),
    .Y(_00803_));
 sky130_vsdinv _16810_ (.A(\cpuregs[1][17] ),
    .Y(_00804_));
 sky130_vsdinv _16811_ (.A(\cpuregs[2][17] ),
    .Y(_00805_));
 sky130_vsdinv _16812_ (.A(\cpuregs[3][17] ),
    .Y(_00806_));
 sky130_vsdinv _16813_ (.A(\cpuregs[4][17] ),
    .Y(_00808_));
 sky130_vsdinv _16814_ (.A(\cpuregs[5][17] ),
    .Y(_00809_));
 sky130_vsdinv _16815_ (.A(\cpuregs[6][17] ),
    .Y(_00810_));
 sky130_vsdinv _16816_ (.A(\cpuregs[7][17] ),
    .Y(_00811_));
 sky130_vsdinv _16817_ (.A(\cpuregs[8][17] ),
    .Y(_00813_));
 sky130_vsdinv _16818_ (.A(\cpuregs[9][17] ),
    .Y(_00814_));
 sky130_vsdinv _16819_ (.A(\cpuregs[10][17] ),
    .Y(_00815_));
 sky130_vsdinv _16820_ (.A(\cpuregs[11][17] ),
    .Y(_00816_));
 sky130_vsdinv _16821_ (.A(\cpuregs[12][17] ),
    .Y(_00818_));
 sky130_vsdinv _16822_ (.A(\cpuregs[13][17] ),
    .Y(_00819_));
 sky130_vsdinv _16823_ (.A(\cpuregs[14][17] ),
    .Y(_00820_));
 sky130_vsdinv _16824_ (.A(\cpuregs[15][17] ),
    .Y(_00821_));
 sky130_vsdinv _16825_ (.A(\cpuregs[16][17] ),
    .Y(_00824_));
 sky130_vsdinv _16826_ (.A(\cpuregs[17][17] ),
    .Y(_00825_));
 sky130_vsdinv _16827_ (.A(\cpuregs[18][17] ),
    .Y(_00826_));
 sky130_vsdinv _16828_ (.A(\cpuregs[19][17] ),
    .Y(_00827_));
 sky130_vsdinv _16829_ (.A(\cpuregs[0][18] ),
    .Y(_00830_));
 sky130_vsdinv _16830_ (.A(\cpuregs[1][18] ),
    .Y(_00831_));
 sky130_vsdinv _16831_ (.A(\cpuregs[2][18] ),
    .Y(_00832_));
 sky130_vsdinv _16832_ (.A(\cpuregs[3][18] ),
    .Y(_00833_));
 sky130_vsdinv _16833_ (.A(\cpuregs[4][18] ),
    .Y(_00835_));
 sky130_vsdinv _16834_ (.A(\cpuregs[5][18] ),
    .Y(_00836_));
 sky130_vsdinv _16835_ (.A(\cpuregs[6][18] ),
    .Y(_00837_));
 sky130_vsdinv _16836_ (.A(\cpuregs[7][18] ),
    .Y(_00838_));
 sky130_vsdinv _16837_ (.A(\cpuregs[8][18] ),
    .Y(_00840_));
 sky130_vsdinv _16838_ (.A(\cpuregs[9][18] ),
    .Y(_00841_));
 sky130_vsdinv _16839_ (.A(\cpuregs[10][18] ),
    .Y(_00842_));
 sky130_vsdinv _16840_ (.A(\cpuregs[11][18] ),
    .Y(_00843_));
 sky130_vsdinv _16841_ (.A(\cpuregs[12][18] ),
    .Y(_00845_));
 sky130_vsdinv _16842_ (.A(\cpuregs[13][18] ),
    .Y(_00846_));
 sky130_vsdinv _16843_ (.A(\cpuregs[14][18] ),
    .Y(_00847_));
 sky130_vsdinv _16844_ (.A(\cpuregs[15][18] ),
    .Y(_00848_));
 sky130_vsdinv _16845_ (.A(\cpuregs[16][18] ),
    .Y(_00851_));
 sky130_vsdinv _16846_ (.A(\cpuregs[17][18] ),
    .Y(_00852_));
 sky130_vsdinv _16847_ (.A(\cpuregs[18][18] ),
    .Y(_00853_));
 sky130_vsdinv _16848_ (.A(\cpuregs[19][18] ),
    .Y(_00854_));
 sky130_vsdinv _16849_ (.A(\cpuregs[0][19] ),
    .Y(_00857_));
 sky130_vsdinv _16850_ (.A(\cpuregs[1][19] ),
    .Y(_00858_));
 sky130_vsdinv _16851_ (.A(\cpuregs[2][19] ),
    .Y(_00859_));
 sky130_vsdinv _16852_ (.A(\cpuregs[3][19] ),
    .Y(_00860_));
 sky130_vsdinv _16853_ (.A(\cpuregs[4][19] ),
    .Y(_00862_));
 sky130_vsdinv _16854_ (.A(\cpuregs[5][19] ),
    .Y(_00863_));
 sky130_vsdinv _16855_ (.A(\cpuregs[6][19] ),
    .Y(_00864_));
 sky130_vsdinv _16856_ (.A(\cpuregs[7][19] ),
    .Y(_00865_));
 sky130_vsdinv _16857_ (.A(\cpuregs[8][19] ),
    .Y(_00867_));
 sky130_vsdinv _16858_ (.A(\cpuregs[9][19] ),
    .Y(_00868_));
 sky130_vsdinv _16859_ (.A(\cpuregs[10][19] ),
    .Y(_00869_));
 sky130_vsdinv _16860_ (.A(\cpuregs[11][19] ),
    .Y(_00870_));
 sky130_vsdinv _16861_ (.A(\cpuregs[12][19] ),
    .Y(_00872_));
 sky130_vsdinv _16862_ (.A(\cpuregs[13][19] ),
    .Y(_00873_));
 sky130_vsdinv _16863_ (.A(\cpuregs[14][19] ),
    .Y(_00874_));
 sky130_vsdinv _16864_ (.A(\cpuregs[15][19] ),
    .Y(_00875_));
 sky130_vsdinv _16865_ (.A(\cpuregs[16][19] ),
    .Y(_00878_));
 sky130_vsdinv _16866_ (.A(\cpuregs[17][19] ),
    .Y(_00879_));
 sky130_vsdinv _16867_ (.A(\cpuregs[18][19] ),
    .Y(_00880_));
 sky130_vsdinv _16868_ (.A(\cpuregs[19][19] ),
    .Y(_00881_));
 sky130_vsdinv _16869_ (.A(\cpuregs[0][20] ),
    .Y(_00884_));
 sky130_vsdinv _16870_ (.A(\cpuregs[1][20] ),
    .Y(_00885_));
 sky130_vsdinv _16871_ (.A(\cpuregs[2][20] ),
    .Y(_00886_));
 sky130_vsdinv _16872_ (.A(\cpuregs[3][20] ),
    .Y(_00887_));
 sky130_vsdinv _16873_ (.A(\cpuregs[4][20] ),
    .Y(_00889_));
 sky130_vsdinv _16874_ (.A(\cpuregs[5][20] ),
    .Y(_00890_));
 sky130_vsdinv _16875_ (.A(\cpuregs[6][20] ),
    .Y(_00891_));
 sky130_vsdinv _16876_ (.A(\cpuregs[7][20] ),
    .Y(_00892_));
 sky130_vsdinv _16877_ (.A(\cpuregs[8][20] ),
    .Y(_00894_));
 sky130_vsdinv _16878_ (.A(\cpuregs[9][20] ),
    .Y(_00895_));
 sky130_vsdinv _16879_ (.A(\cpuregs[10][20] ),
    .Y(_00896_));
 sky130_vsdinv _16880_ (.A(\cpuregs[11][20] ),
    .Y(_00897_));
 sky130_vsdinv _16881_ (.A(\cpuregs[12][20] ),
    .Y(_00899_));
 sky130_vsdinv _16882_ (.A(\cpuregs[13][20] ),
    .Y(_00900_));
 sky130_vsdinv _16883_ (.A(\cpuregs[14][20] ),
    .Y(_00901_));
 sky130_vsdinv _16884_ (.A(\cpuregs[15][20] ),
    .Y(_00902_));
 sky130_vsdinv _16885_ (.A(\cpuregs[16][20] ),
    .Y(_00905_));
 sky130_vsdinv _16886_ (.A(\cpuregs[17][20] ),
    .Y(_00906_));
 sky130_vsdinv _16887_ (.A(\cpuregs[18][20] ),
    .Y(_00907_));
 sky130_vsdinv _16888_ (.A(\cpuregs[19][20] ),
    .Y(_00908_));
 sky130_vsdinv _16889_ (.A(\cpuregs[0][21] ),
    .Y(_00911_));
 sky130_vsdinv _16890_ (.A(\cpuregs[1][21] ),
    .Y(_00912_));
 sky130_vsdinv _16891_ (.A(\cpuregs[2][21] ),
    .Y(_00913_));
 sky130_vsdinv _16892_ (.A(\cpuregs[3][21] ),
    .Y(_00914_));
 sky130_vsdinv _16893_ (.A(\cpuregs[4][21] ),
    .Y(_00916_));
 sky130_vsdinv _16894_ (.A(\cpuregs[5][21] ),
    .Y(_00917_));
 sky130_vsdinv _16895_ (.A(\cpuregs[6][21] ),
    .Y(_00918_));
 sky130_vsdinv _16896_ (.A(\cpuregs[7][21] ),
    .Y(_00919_));
 sky130_vsdinv _16897_ (.A(\cpuregs[8][21] ),
    .Y(_00921_));
 sky130_vsdinv _16898_ (.A(\cpuregs[9][21] ),
    .Y(_00922_));
 sky130_vsdinv _16899_ (.A(\cpuregs[10][21] ),
    .Y(_00923_));
 sky130_vsdinv _16900_ (.A(\cpuregs[11][21] ),
    .Y(_00924_));
 sky130_vsdinv _16901_ (.A(\cpuregs[12][21] ),
    .Y(_00926_));
 sky130_vsdinv _16902_ (.A(\cpuregs[13][21] ),
    .Y(_00927_));
 sky130_vsdinv _16903_ (.A(\cpuregs[14][21] ),
    .Y(_00928_));
 sky130_vsdinv _16904_ (.A(\cpuregs[15][21] ),
    .Y(_00929_));
 sky130_vsdinv _16905_ (.A(\cpuregs[16][21] ),
    .Y(_00932_));
 sky130_vsdinv _16906_ (.A(\cpuregs[17][21] ),
    .Y(_00933_));
 sky130_vsdinv _16907_ (.A(\cpuregs[18][21] ),
    .Y(_00934_));
 sky130_vsdinv _16908_ (.A(\cpuregs[19][21] ),
    .Y(_00935_));
 sky130_vsdinv _16909_ (.A(\cpuregs[0][22] ),
    .Y(_00938_));
 sky130_vsdinv _16910_ (.A(\cpuregs[1][22] ),
    .Y(_00939_));
 sky130_vsdinv _16911_ (.A(\cpuregs[2][22] ),
    .Y(_00940_));
 sky130_vsdinv _16912_ (.A(\cpuregs[3][22] ),
    .Y(_00941_));
 sky130_vsdinv _16913_ (.A(\cpuregs[4][22] ),
    .Y(_00943_));
 sky130_vsdinv _16914_ (.A(\cpuregs[5][22] ),
    .Y(_00944_));
 sky130_vsdinv _16915_ (.A(\cpuregs[6][22] ),
    .Y(_00945_));
 sky130_vsdinv _16916_ (.A(\cpuregs[7][22] ),
    .Y(_00946_));
 sky130_fd_sc_hd__o32a_2 _16917_ (.A1(_11779_),
    .A2(_11807_),
    .A3(_10809_),
    .B1(_11786_),
    .B2(_10812_),
    .X(_12370_));
 sky130_fd_sc_hd__or2_2 _16918_ (.A(_00296_),
    .B(_12370_),
    .X(_12371_));
 sky130_fd_sc_hd__o221ai_2 _16919_ (.A1(_10689_),
    .A2(_00322_),
    .B1(_12209_),
    .B2(_12363_),
    .C1(_12371_),
    .Y(_00045_));
 sky130_vsdinv _16920_ (.A(\cpuregs[8][22] ),
    .Y(_00948_));
 sky130_vsdinv _16921_ (.A(\cpuregs[9][22] ),
    .Y(_00949_));
 sky130_vsdinv _16922_ (.A(\cpuregs[10][22] ),
    .Y(_00950_));
 sky130_vsdinv _16923_ (.A(\cpuregs[11][22] ),
    .Y(_00951_));
 sky130_vsdinv _16924_ (.A(\cpuregs[12][22] ),
    .Y(_00953_));
 sky130_vsdinv _16925_ (.A(\cpuregs[13][22] ),
    .Y(_00954_));
 sky130_vsdinv _16926_ (.A(\cpuregs[14][22] ),
    .Y(_00955_));
 sky130_vsdinv _16927_ (.A(\cpuregs[15][22] ),
    .Y(_00956_));
 sky130_vsdinv _16928_ (.A(\cpuregs[16][22] ),
    .Y(_00959_));
 sky130_vsdinv _16929_ (.A(\cpuregs[17][22] ),
    .Y(_00960_));
 sky130_vsdinv _16930_ (.A(\cpuregs[18][22] ),
    .Y(_00961_));
 sky130_vsdinv _16931_ (.A(\cpuregs[19][22] ),
    .Y(_00962_));
 sky130_vsdinv _16932_ (.A(\cpuregs[0][23] ),
    .Y(_00965_));
 sky130_vsdinv _16933_ (.A(\cpuregs[1][23] ),
    .Y(_00966_));
 sky130_vsdinv _16934_ (.A(\cpuregs[2][23] ),
    .Y(_00967_));
 sky130_vsdinv _16935_ (.A(\cpuregs[3][23] ),
    .Y(_00968_));
 sky130_vsdinv _16936_ (.A(\cpuregs[4][23] ),
    .Y(_00970_));
 sky130_vsdinv _16937_ (.A(\cpuregs[5][23] ),
    .Y(_00971_));
 sky130_vsdinv _16938_ (.A(\cpuregs[6][23] ),
    .Y(_00972_));
 sky130_vsdinv _16939_ (.A(\cpuregs[7][23] ),
    .Y(_00973_));
 sky130_vsdinv _16940_ (.A(\cpuregs[8][23] ),
    .Y(_00975_));
 sky130_vsdinv _16941_ (.A(\cpuregs[9][23] ),
    .Y(_00976_));
 sky130_vsdinv _16942_ (.A(\cpuregs[10][23] ),
    .Y(_00977_));
 sky130_vsdinv _16943_ (.A(\cpuregs[11][23] ),
    .Y(_00978_));
 sky130_vsdinv _16944_ (.A(\cpuregs[12][23] ),
    .Y(_00980_));
 sky130_vsdinv _16945_ (.A(\cpuregs[13][23] ),
    .Y(_00981_));
 sky130_vsdinv _16946_ (.A(\cpuregs[14][23] ),
    .Y(_00982_));
 sky130_vsdinv _16947_ (.A(\cpuregs[15][23] ),
    .Y(_00983_));
 sky130_vsdinv _16948_ (.A(\cpuregs[16][23] ),
    .Y(_00986_));
 sky130_vsdinv _16949_ (.A(\cpuregs[17][23] ),
    .Y(_00987_));
 sky130_vsdinv _16950_ (.A(\cpuregs[18][23] ),
    .Y(_00988_));
 sky130_vsdinv _16951_ (.A(\cpuregs[19][23] ),
    .Y(_00989_));
 sky130_vsdinv _16952_ (.A(\cpuregs[0][24] ),
    .Y(_00992_));
 sky130_vsdinv _16953_ (.A(\cpuregs[1][24] ),
    .Y(_00993_));
 sky130_vsdinv _16954_ (.A(\cpuregs[2][24] ),
    .Y(_00994_));
 sky130_vsdinv _16955_ (.A(\cpuregs[3][24] ),
    .Y(_00995_));
 sky130_vsdinv _16956_ (.A(\cpuregs[4][24] ),
    .Y(_00997_));
 sky130_vsdinv _16957_ (.A(\cpuregs[5][24] ),
    .Y(_00998_));
 sky130_vsdinv _16958_ (.A(\cpuregs[6][24] ),
    .Y(_00999_));
 sky130_vsdinv _16959_ (.A(\cpuregs[7][24] ),
    .Y(_01000_));
 sky130_vsdinv _16960_ (.A(\cpuregs[8][24] ),
    .Y(_01002_));
 sky130_vsdinv _16961_ (.A(\cpuregs[9][24] ),
    .Y(_01003_));
 sky130_vsdinv _16962_ (.A(\cpuregs[10][24] ),
    .Y(_01004_));
 sky130_vsdinv _16963_ (.A(\cpuregs[11][24] ),
    .Y(_01005_));
 sky130_vsdinv _16964_ (.A(\cpuregs[12][24] ),
    .Y(_01007_));
 sky130_vsdinv _16965_ (.A(\cpuregs[13][24] ),
    .Y(_01008_));
 sky130_vsdinv _16966_ (.A(\cpuregs[14][24] ),
    .Y(_01009_));
 sky130_vsdinv _16967_ (.A(\cpuregs[15][24] ),
    .Y(_01010_));
 sky130_vsdinv _16968_ (.A(\cpuregs[16][24] ),
    .Y(_01013_));
 sky130_vsdinv _16969_ (.A(\cpuregs[17][24] ),
    .Y(_01014_));
 sky130_vsdinv _16970_ (.A(\cpuregs[18][24] ),
    .Y(_01015_));
 sky130_vsdinv _16971_ (.A(\cpuregs[19][24] ),
    .Y(_01016_));
 sky130_vsdinv _16972_ (.A(\cpuregs[0][25] ),
    .Y(_01019_));
 sky130_vsdinv _16973_ (.A(\cpuregs[1][25] ),
    .Y(_01020_));
 sky130_vsdinv _16974_ (.A(\cpuregs[2][25] ),
    .Y(_01021_));
 sky130_vsdinv _16975_ (.A(\cpuregs[3][25] ),
    .Y(_01022_));
 sky130_vsdinv _16976_ (.A(\cpuregs[4][25] ),
    .Y(_01024_));
 sky130_vsdinv _16977_ (.A(\cpuregs[5][25] ),
    .Y(_01025_));
 sky130_vsdinv _16978_ (.A(\cpuregs[6][25] ),
    .Y(_01026_));
 sky130_vsdinv _16979_ (.A(\cpuregs[7][25] ),
    .Y(_01027_));
 sky130_fd_sc_hd__nor2_2 _16980_ (.A(\mem_state[1] ),
    .B(_10449_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_2 _16981_ (.A(_10480_),
    .B(_00289_),
    .Y(_00298_));
 sky130_vsdinv _16982_ (.A(\cpuregs[8][25] ),
    .Y(_01029_));
 sky130_vsdinv _16983_ (.A(\cpuregs[9][25] ),
    .Y(_01030_));
 sky130_vsdinv _16984_ (.A(\cpuregs[10][25] ),
    .Y(_01031_));
 sky130_vsdinv _16985_ (.A(\cpuregs[11][25] ),
    .Y(_01032_));
 sky130_vsdinv _16986_ (.A(\cpuregs[12][25] ),
    .Y(_01034_));
 sky130_vsdinv _16987_ (.A(\cpuregs[13][25] ),
    .Y(_01035_));
 sky130_vsdinv _16988_ (.A(\cpuregs[14][25] ),
    .Y(_01036_));
 sky130_vsdinv _16989_ (.A(\cpuregs[15][25] ),
    .Y(_01037_));
 sky130_vsdinv _16990_ (.A(\cpuregs[16][25] ),
    .Y(_01040_));
 sky130_vsdinv _16991_ (.A(\cpuregs[17][25] ),
    .Y(_01041_));
 sky130_vsdinv _16992_ (.A(\cpuregs[18][25] ),
    .Y(_01042_));
 sky130_vsdinv _16993_ (.A(\cpuregs[19][25] ),
    .Y(_01043_));
 sky130_vsdinv _16994_ (.A(\cpuregs[0][26] ),
    .Y(_01046_));
 sky130_vsdinv _16995_ (.A(\cpuregs[1][26] ),
    .Y(_01047_));
 sky130_vsdinv _16996_ (.A(\cpuregs[2][26] ),
    .Y(_01048_));
 sky130_vsdinv _16997_ (.A(\cpuregs[3][26] ),
    .Y(_01049_));
 sky130_vsdinv _16998_ (.A(\cpuregs[4][26] ),
    .Y(_01051_));
 sky130_vsdinv _16999_ (.A(\cpuregs[5][26] ),
    .Y(_01052_));
 sky130_vsdinv _17000_ (.A(\cpuregs[6][26] ),
    .Y(_01053_));
 sky130_vsdinv _17001_ (.A(\cpuregs[7][26] ),
    .Y(_01054_));
 sky130_vsdinv _17002_ (.A(\cpuregs[8][26] ),
    .Y(_01056_));
 sky130_vsdinv _17003_ (.A(\cpuregs[9][26] ),
    .Y(_01057_));
 sky130_vsdinv _17004_ (.A(\cpuregs[10][26] ),
    .Y(_01058_));
 sky130_vsdinv _17005_ (.A(\cpuregs[11][26] ),
    .Y(_01059_));
 sky130_vsdinv _17006_ (.A(\cpuregs[12][26] ),
    .Y(_01061_));
 sky130_vsdinv _17007_ (.A(\cpuregs[13][26] ),
    .Y(_01062_));
 sky130_vsdinv _17008_ (.A(\cpuregs[14][26] ),
    .Y(_01063_));
 sky130_vsdinv _17009_ (.A(\cpuregs[15][26] ),
    .Y(_01064_));
 sky130_vsdinv _17010_ (.A(\cpuregs[16][26] ),
    .Y(_01067_));
 sky130_vsdinv _17011_ (.A(\cpuregs[17][26] ),
    .Y(_01068_));
 sky130_vsdinv _17012_ (.A(\cpuregs[18][26] ),
    .Y(_01069_));
 sky130_vsdinv _17013_ (.A(\cpuregs[19][26] ),
    .Y(_01070_));
 sky130_vsdinv _17014_ (.A(\mem_wordsize[1] ),
    .Y(_12372_));
 sky130_fd_sc_hd__buf_1 _17015_ (.A(_12372_),
    .X(_12373_));
 sky130_fd_sc_hd__o211a_2 _17016_ (.A1(instr_lbu),
    .A2(instr_lb),
    .B1(_10456_),
    .C1(_10457_),
    .X(_12374_));
 sky130_fd_sc_hd__a31oi_2 _17017_ (.A1(_00291_),
    .A2(instr_sb),
    .A3(\cpu_state[5] ),
    .B1(_12374_),
    .Y(_12375_));
 sky130_fd_sc_hd__o22ai_2 _17018_ (.A1(_12373_),
    .A2(_12363_),
    .B1(_12259_),
    .B2(_12375_),
    .Y(_00046_));
 sky130_vsdinv _17019_ (.A(\cpuregs[0][27] ),
    .Y(_01073_));
 sky130_vsdinv _17020_ (.A(\cpuregs[1][27] ),
    .Y(_01074_));
 sky130_vsdinv _17021_ (.A(\cpuregs[2][27] ),
    .Y(_01075_));
 sky130_vsdinv _17022_ (.A(\cpuregs[3][27] ),
    .Y(_01076_));
 sky130_vsdinv _17023_ (.A(\cpuregs[4][27] ),
    .Y(_01078_));
 sky130_vsdinv _17024_ (.A(\cpuregs[5][27] ),
    .Y(_01079_));
 sky130_vsdinv _17025_ (.A(\cpuregs[6][27] ),
    .Y(_01080_));
 sky130_vsdinv _17026_ (.A(\cpuregs[7][27] ),
    .Y(_01081_));
 sky130_vsdinv _17027_ (.A(\cpuregs[8][27] ),
    .Y(_01083_));
 sky130_vsdinv _17028_ (.A(\cpuregs[9][27] ),
    .Y(_01084_));
 sky130_vsdinv _17029_ (.A(\cpuregs[10][27] ),
    .Y(_01085_));
 sky130_vsdinv _17030_ (.A(\cpuregs[11][27] ),
    .Y(_01086_));
 sky130_vsdinv _17031_ (.A(\cpuregs[12][27] ),
    .Y(_01088_));
 sky130_vsdinv _17032_ (.A(\cpuregs[13][27] ),
    .Y(_01089_));
 sky130_vsdinv _17033_ (.A(\cpuregs[14][27] ),
    .Y(_01090_));
 sky130_vsdinv _17034_ (.A(\cpuregs[15][27] ),
    .Y(_01091_));
 sky130_vsdinv _17035_ (.A(\cpuregs[16][27] ),
    .Y(_01094_));
 sky130_vsdinv _17036_ (.A(\cpuregs[17][27] ),
    .Y(_01095_));
 sky130_vsdinv _17037_ (.A(\cpuregs[18][27] ),
    .Y(_01096_));
 sky130_vsdinv _17038_ (.A(\cpuregs[19][27] ),
    .Y(_01097_));
 sky130_vsdinv _17039_ (.A(\cpuregs[0][28] ),
    .Y(_01100_));
 sky130_vsdinv _17040_ (.A(\cpuregs[1][28] ),
    .Y(_01101_));
 sky130_vsdinv _17041_ (.A(\cpuregs[2][28] ),
    .Y(_01102_));
 sky130_vsdinv _17042_ (.A(\cpuregs[3][28] ),
    .Y(_01103_));
 sky130_vsdinv _17043_ (.A(\cpuregs[4][28] ),
    .Y(_01105_));
 sky130_vsdinv _17044_ (.A(\cpuregs[5][28] ),
    .Y(_01106_));
 sky130_vsdinv _17045_ (.A(\cpuregs[6][28] ),
    .Y(_01107_));
 sky130_vsdinv _17046_ (.A(\cpuregs[7][28] ),
    .Y(_01108_));
 sky130_vsdinv _17047_ (.A(\cpuregs[8][28] ),
    .Y(_01110_));
 sky130_vsdinv _17048_ (.A(\cpuregs[9][28] ),
    .Y(_01111_));
 sky130_vsdinv _17049_ (.A(\cpuregs[10][28] ),
    .Y(_01112_));
 sky130_vsdinv _17050_ (.A(\cpuregs[11][28] ),
    .Y(_01113_));
 sky130_vsdinv _17051_ (.A(\cpuregs[12][28] ),
    .Y(_01115_));
 sky130_vsdinv _17052_ (.A(\cpuregs[13][28] ),
    .Y(_01116_));
 sky130_vsdinv _17053_ (.A(\cpuregs[14][28] ),
    .Y(_01117_));
 sky130_vsdinv _17054_ (.A(\cpuregs[15][28] ),
    .Y(_01118_));
 sky130_vsdinv _17055_ (.A(\cpuregs[16][28] ),
    .Y(_01121_));
 sky130_vsdinv _17056_ (.A(\cpuregs[17][28] ),
    .Y(_01122_));
 sky130_vsdinv _17057_ (.A(\cpuregs[18][28] ),
    .Y(_01123_));
 sky130_vsdinv _17058_ (.A(\cpuregs[19][28] ),
    .Y(_01124_));
 sky130_vsdinv _17059_ (.A(\cpuregs[0][29] ),
    .Y(_01127_));
 sky130_vsdinv _17060_ (.A(\cpuregs[1][29] ),
    .Y(_01128_));
 sky130_vsdinv _17061_ (.A(\cpuregs[2][29] ),
    .Y(_01129_));
 sky130_vsdinv _17062_ (.A(\cpuregs[3][29] ),
    .Y(_01130_));
 sky130_vsdinv _17063_ (.A(\cpuregs[4][29] ),
    .Y(_01132_));
 sky130_vsdinv _17064_ (.A(\cpuregs[5][29] ),
    .Y(_01133_));
 sky130_vsdinv _17065_ (.A(\cpuregs[6][29] ),
    .Y(_01134_));
 sky130_vsdinv _17066_ (.A(\cpuregs[7][29] ),
    .Y(_01135_));
 sky130_vsdinv _17067_ (.A(\cpuregs[8][29] ),
    .Y(_01137_));
 sky130_vsdinv _17068_ (.A(\cpuregs[9][29] ),
    .Y(_01138_));
 sky130_vsdinv _17069_ (.A(\cpuregs[10][29] ),
    .Y(_01139_));
 sky130_vsdinv _17070_ (.A(\cpuregs[11][29] ),
    .Y(_01140_));
 sky130_vsdinv _17071_ (.A(\cpuregs[12][29] ),
    .Y(_01142_));
 sky130_vsdinv _17072_ (.A(\cpuregs[13][29] ),
    .Y(_01143_));
 sky130_fd_sc_hd__buf_1 _17073_ (.A(_10473_),
    .X(_12376_));
 sky130_fd_sc_hd__and2_2 _17074_ (.A(_12376_),
    .B(_00294_),
    .X(_00295_));
 sky130_vsdinv _17075_ (.A(\cpuregs[14][29] ),
    .Y(_01144_));
 sky130_vsdinv _17076_ (.A(\cpuregs[15][29] ),
    .Y(_01145_));
 sky130_vsdinv _17077_ (.A(\cpuregs[16][29] ),
    .Y(_01148_));
 sky130_vsdinv _17078_ (.A(\cpuregs[17][29] ),
    .Y(_01149_));
 sky130_vsdinv _17079_ (.A(\cpuregs[18][29] ),
    .Y(_01150_));
 sky130_vsdinv _17080_ (.A(\cpuregs[19][29] ),
    .Y(_01151_));
 sky130_vsdinv _17081_ (.A(\cpuregs[0][30] ),
    .Y(_01154_));
 sky130_vsdinv _17082_ (.A(\cpuregs[1][30] ),
    .Y(_01155_));
 sky130_vsdinv _17083_ (.A(\cpuregs[2][30] ),
    .Y(_01156_));
 sky130_vsdinv _17084_ (.A(\cpuregs[3][30] ),
    .Y(_01157_));
 sky130_vsdinv _17085_ (.A(\cpuregs[4][30] ),
    .Y(_01159_));
 sky130_vsdinv _17086_ (.A(\cpuregs[5][30] ),
    .Y(_01160_));
 sky130_vsdinv _17087_ (.A(\cpuregs[6][30] ),
    .Y(_01161_));
 sky130_vsdinv _17088_ (.A(\cpuregs[7][30] ),
    .Y(_01162_));
 sky130_vsdinv _17089_ (.A(\cpuregs[8][30] ),
    .Y(_01164_));
 sky130_vsdinv _17090_ (.A(\cpuregs[9][30] ),
    .Y(_01165_));
 sky130_vsdinv _17091_ (.A(\cpuregs[10][30] ),
    .Y(_01166_));
 sky130_vsdinv _17092_ (.A(\cpuregs[11][30] ),
    .Y(_01167_));
 sky130_vsdinv _17093_ (.A(\cpuregs[12][30] ),
    .Y(_01169_));
 sky130_vsdinv _17094_ (.A(\cpuregs[13][30] ),
    .Y(_01170_));
 sky130_vsdinv _17095_ (.A(\cpuregs[14][30] ),
    .Y(_01171_));
 sky130_vsdinv _17096_ (.A(\cpuregs[15][30] ),
    .Y(_01172_));
 sky130_vsdinv _17097_ (.A(\cpuregs[16][30] ),
    .Y(_01175_));
 sky130_vsdinv _17098_ (.A(\cpuregs[17][30] ),
    .Y(_01176_));
 sky130_vsdinv _17099_ (.A(\cpuregs[18][30] ),
    .Y(_01177_));
 sky130_vsdinv _17100_ (.A(\cpuregs[19][30] ),
    .Y(_01178_));
 sky130_vsdinv _17101_ (.A(\cpuregs[0][31] ),
    .Y(_01181_));
 sky130_vsdinv _17102_ (.A(\cpuregs[1][31] ),
    .Y(_01182_));
 sky130_vsdinv _17103_ (.A(\cpuregs[2][31] ),
    .Y(_01183_));
 sky130_vsdinv _17104_ (.A(\cpuregs[3][31] ),
    .Y(_01184_));
 sky130_vsdinv _17105_ (.A(\cpuregs[4][31] ),
    .Y(_01186_));
 sky130_vsdinv _17106_ (.A(\cpuregs[5][31] ),
    .Y(_01187_));
 sky130_vsdinv _17107_ (.A(\cpuregs[6][31] ),
    .Y(_01188_));
 sky130_vsdinv _17108_ (.A(\cpuregs[7][31] ),
    .Y(_01189_));
 sky130_vsdinv _17109_ (.A(\cpuregs[8][31] ),
    .Y(_01191_));
 sky130_vsdinv _17110_ (.A(\cpuregs[9][31] ),
    .Y(_01192_));
 sky130_vsdinv _17111_ (.A(\cpuregs[10][31] ),
    .Y(_01193_));
 sky130_vsdinv _17112_ (.A(\cpuregs[11][31] ),
    .Y(_01194_));
 sky130_vsdinv _17113_ (.A(\cpuregs[12][31] ),
    .Y(_01196_));
 sky130_vsdinv _17114_ (.A(\cpuregs[13][31] ),
    .Y(_01197_));
 sky130_vsdinv _17115_ (.A(\cpuregs[14][31] ),
    .Y(_01198_));
 sky130_vsdinv _17116_ (.A(\cpuregs[15][31] ),
    .Y(_01199_));
 sky130_vsdinv _17117_ (.A(\cpuregs[16][31] ),
    .Y(_01202_));
 sky130_vsdinv _17118_ (.A(\cpuregs[17][31] ),
    .Y(_01203_));
 sky130_vsdinv _17119_ (.A(\cpuregs[18][31] ),
    .Y(_01204_));
 sky130_vsdinv _17120_ (.A(\cpuregs[19][31] ),
    .Y(_01205_));
 sky130_vsdinv _17121_ (.A(\timer[26] ),
    .Y(_12377_));
 sky130_vsdinv _17122_ (.A(\timer[18] ),
    .Y(_12378_));
 sky130_fd_sc_hd__or2_2 _17123_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .X(_12379_));
 sky130_fd_sc_hd__or2_2 _17124_ (.A(\timer[2] ),
    .B(_12379_),
    .X(_12380_));
 sky130_fd_sc_hd__or2_2 _17125_ (.A(\timer[3] ),
    .B(_12380_),
    .X(_12381_));
 sky130_fd_sc_hd__or3_2 _17126_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .C(_12381_),
    .X(_12382_));
 sky130_fd_sc_hd__or2_2 _17127_ (.A(\timer[6] ),
    .B(_12382_),
    .X(_12383_));
 sky130_fd_sc_hd__or2_2 _17128_ (.A(\timer[7] ),
    .B(_12383_),
    .X(_12384_));
 sky130_fd_sc_hd__or2_2 _17129_ (.A(\timer[8] ),
    .B(_12384_),
    .X(_12385_));
 sky130_fd_sc_hd__or2_2 _17130_ (.A(\timer[9] ),
    .B(_12385_),
    .X(_12386_));
 sky130_fd_sc_hd__or2_2 _17131_ (.A(\timer[10] ),
    .B(_12386_),
    .X(_12387_));
 sky130_fd_sc_hd__or2_2 _17132_ (.A(\timer[11] ),
    .B(_12387_),
    .X(_12388_));
 sky130_fd_sc_hd__or2_2 _17133_ (.A(\timer[12] ),
    .B(_12388_),
    .X(_12389_));
 sky130_fd_sc_hd__or2_2 _17134_ (.A(\timer[13] ),
    .B(_12389_),
    .X(_12390_));
 sky130_fd_sc_hd__or2_2 _17135_ (.A(\timer[14] ),
    .B(_12390_),
    .X(_12391_));
 sky130_fd_sc_hd__or2_2 _17136_ (.A(\timer[15] ),
    .B(_12391_),
    .X(_12392_));
 sky130_fd_sc_hd__or2_2 _17137_ (.A(\timer[16] ),
    .B(_12392_),
    .X(_12393_));
 sky130_fd_sc_hd__nor2_2 _17138_ (.A(\timer[17] ),
    .B(_12393_),
    .Y(_12394_));
 sky130_fd_sc_hd__nand2_2 _17139_ (.A(_12378_),
    .B(_12394_),
    .Y(_12395_));
 sky130_fd_sc_hd__or2_2 _17140_ (.A(\timer[19] ),
    .B(_12395_),
    .X(_12396_));
 sky130_fd_sc_hd__or2_2 _17141_ (.A(\timer[20] ),
    .B(_12396_),
    .X(_12397_));
 sky130_fd_sc_hd__or2_2 _17142_ (.A(\timer[21] ),
    .B(_12397_),
    .X(_12398_));
 sky130_fd_sc_hd__or2_2 _17143_ (.A(\timer[22] ),
    .B(_12398_),
    .X(_12399_));
 sky130_fd_sc_hd__or2_2 _17144_ (.A(\timer[23] ),
    .B(_12399_),
    .X(_12400_));
 sky130_fd_sc_hd__or2_2 _17145_ (.A(\timer[24] ),
    .B(_12400_),
    .X(_12401_));
 sky130_fd_sc_hd__nor2_2 _17146_ (.A(\timer[25] ),
    .B(_12401_),
    .Y(_12402_));
 sky130_fd_sc_hd__nand2_2 _17147_ (.A(_12377_),
    .B(_12402_),
    .Y(_12403_));
 sky130_fd_sc_hd__or2_2 _17148_ (.A(\timer[27] ),
    .B(_12403_),
    .X(_12404_));
 sky130_fd_sc_hd__or2_2 _17149_ (.A(\timer[28] ),
    .B(_12404_),
    .X(_12405_));
 sky130_fd_sc_hd__or2_2 _17150_ (.A(\timer[29] ),
    .B(_12405_),
    .X(_12406_));
 sky130_fd_sc_hd__or2_2 _17151_ (.A(\timer[30] ),
    .B(_12406_),
    .X(_12407_));
 sky130_fd_sc_hd__nor2_2 _17152_ (.A(\timer[31] ),
    .B(_12407_),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_2 _17153_ (.A(\timer[0] ),
    .B(_01208_),
    .Y(_01209_));
 sky130_vsdinv _17154_ (.A(\timer[1] ),
    .Y(_12408_));
 sky130_vsdinv _17155_ (.A(\timer[0] ),
    .Y(_12409_));
 sky130_fd_sc_hd__o21ai_2 _17156_ (.A1(_12408_),
    .A2(_12409_),
    .B1(_12379_),
    .Y(_01211_));
 sky130_fd_sc_hd__a21bo_2 _17157_ (.A1(\timer[2] ),
    .A2(_12379_),
    .B1_N(_12380_),
    .X(_01214_));
 sky130_fd_sc_hd__a21bo_2 _17158_ (.A1(\timer[3] ),
    .A2(_12380_),
    .B1_N(_12381_),
    .X(_01217_));
 sky130_fd_sc_hd__nor2_2 _17159_ (.A(\timer[4] ),
    .B(_12381_),
    .Y(_12410_));
 sky130_fd_sc_hd__a21o_2 _17160_ (.A1(\timer[4] ),
    .A2(_12381_),
    .B1(_12410_),
    .X(_01220_));
 sky130_vsdinv _17161_ (.A(\timer[5] ),
    .Y(_12411_));
 sky130_fd_sc_hd__o21ai_2 _17162_ (.A1(_12411_),
    .A2(_12410_),
    .B1(_12382_),
    .Y(_01223_));
 sky130_vsdinv _17163_ (.A(_12383_),
    .Y(_12412_));
 sky130_fd_sc_hd__a21o_2 _17164_ (.A1(\timer[6] ),
    .A2(_12382_),
    .B1(_12412_),
    .X(_01226_));
 sky130_vsdinv _17165_ (.A(\timer[7] ),
    .Y(_12413_));
 sky130_fd_sc_hd__o21ai_2 _17166_ (.A1(_12413_),
    .A2(_12412_),
    .B1(_12384_),
    .Y(_01229_));
 sky130_vsdinv _17167_ (.A(_12385_),
    .Y(_12414_));
 sky130_fd_sc_hd__a21o_2 _17168_ (.A1(\timer[8] ),
    .A2(_12384_),
    .B1(_12414_),
    .X(_01232_));
 sky130_vsdinv _17169_ (.A(\timer[9] ),
    .Y(_12415_));
 sky130_fd_sc_hd__o21ai_2 _17170_ (.A1(_12415_),
    .A2(_12414_),
    .B1(_12386_),
    .Y(_01235_));
 sky130_vsdinv _17171_ (.A(_12387_),
    .Y(_12416_));
 sky130_fd_sc_hd__a21o_2 _17172_ (.A1(\timer[10] ),
    .A2(_12386_),
    .B1(_12416_),
    .X(_01238_));
 sky130_vsdinv _17173_ (.A(\timer[11] ),
    .Y(_12417_));
 sky130_fd_sc_hd__o21ai_2 _17174_ (.A1(_12417_),
    .A2(_12416_),
    .B1(_12388_),
    .Y(_01241_));
 sky130_vsdinv _17175_ (.A(_12389_),
    .Y(_12418_));
 sky130_fd_sc_hd__a21o_2 _17176_ (.A1(\timer[12] ),
    .A2(_12388_),
    .B1(_12418_),
    .X(_01244_));
 sky130_vsdinv _17177_ (.A(\timer[13] ),
    .Y(_12419_));
 sky130_fd_sc_hd__o21ai_2 _17178_ (.A1(_12419_),
    .A2(_12418_),
    .B1(_12390_),
    .Y(_01247_));
 sky130_vsdinv _17179_ (.A(_12391_),
    .Y(_12420_));
 sky130_fd_sc_hd__a21o_2 _17180_ (.A1(\timer[14] ),
    .A2(_12390_),
    .B1(_12420_),
    .X(_01250_));
 sky130_vsdinv _17181_ (.A(\timer[15] ),
    .Y(_12421_));
 sky130_fd_sc_hd__o21ai_2 _17182_ (.A1(_12421_),
    .A2(_12420_),
    .B1(_12392_),
    .Y(_01253_));
 sky130_fd_sc_hd__a21bo_2 _17183_ (.A1(\timer[16] ),
    .A2(_12392_),
    .B1_N(_12393_),
    .X(_01256_));
 sky130_fd_sc_hd__a21o_2 _17184_ (.A1(\timer[17] ),
    .A2(_12393_),
    .B1(_12394_),
    .X(_01259_));
 sky130_fd_sc_hd__o21ai_2 _17185_ (.A1(_12378_),
    .A2(_12394_),
    .B1(_12395_),
    .Y(_01262_));
 sky130_vsdinv _17186_ (.A(_12396_),
    .Y(_12422_));
 sky130_fd_sc_hd__a21o_2 _17187_ (.A1(\timer[19] ),
    .A2(_12395_),
    .B1(_12422_),
    .X(_01265_));
 sky130_vsdinv _17188_ (.A(\timer[20] ),
    .Y(_12423_));
 sky130_fd_sc_hd__o21ai_2 _17189_ (.A1(_12423_),
    .A2(_12422_),
    .B1(_12397_),
    .Y(_01268_));
 sky130_vsdinv _17190_ (.A(_12398_),
    .Y(_12424_));
 sky130_fd_sc_hd__a21o_2 _17191_ (.A1(\timer[21] ),
    .A2(_12397_),
    .B1(_12424_),
    .X(_01271_));
 sky130_vsdinv _17192_ (.A(\timer[22] ),
    .Y(_12425_));
 sky130_fd_sc_hd__o21ai_2 _17193_ (.A1(_12425_),
    .A2(_12424_),
    .B1(_12399_),
    .Y(_01274_));
 sky130_vsdinv _17194_ (.A(_12400_),
    .Y(_12426_));
 sky130_fd_sc_hd__a21o_2 _17195_ (.A1(\timer[23] ),
    .A2(_12399_),
    .B1(_12426_),
    .X(_01277_));
 sky130_vsdinv _17196_ (.A(\timer[24] ),
    .Y(_12427_));
 sky130_fd_sc_hd__o21ai_2 _17197_ (.A1(_12427_),
    .A2(_12426_),
    .B1(_12401_),
    .Y(_01280_));
 sky130_fd_sc_hd__a21o_2 _17198_ (.A1(\timer[25] ),
    .A2(_12401_),
    .B1(_12402_),
    .X(_01283_));
 sky130_fd_sc_hd__o21ai_2 _17199_ (.A1(_12377_),
    .A2(_12402_),
    .B1(_12403_),
    .Y(_01286_));
 sky130_vsdinv _17200_ (.A(_12404_),
    .Y(_12428_));
 sky130_fd_sc_hd__a21o_2 _17201_ (.A1(\timer[27] ),
    .A2(_12403_),
    .B1(_12428_),
    .X(_01289_));
 sky130_vsdinv _17202_ (.A(\timer[28] ),
    .Y(_12429_));
 sky130_fd_sc_hd__o21ai_2 _17203_ (.A1(_12429_),
    .A2(_12428_),
    .B1(_12405_),
    .Y(_01292_));
 sky130_vsdinv _17204_ (.A(_12406_),
    .Y(_12430_));
 sky130_fd_sc_hd__a21o_2 _17205_ (.A1(\timer[29] ),
    .A2(_12405_),
    .B1(_12430_),
    .X(_01295_));
 sky130_vsdinv _17206_ (.A(\timer[30] ),
    .Y(_12431_));
 sky130_fd_sc_hd__o21ai_2 _17207_ (.A1(_12431_),
    .A2(_12430_),
    .B1(_12407_),
    .Y(_01298_));
 sky130_fd_sc_hd__a21o_2 _17208_ (.A1(\timer[31] ),
    .A2(_12407_),
    .B1(_01208_),
    .X(_01301_));
 sky130_fd_sc_hd__nor2_2 _17209_ (.A(_11700_),
    .B(_12084_),
    .Y(_01315_));
 sky130_fd_sc_hd__nor2_2 _17210_ (.A(_11700_),
    .B(_12091_),
    .Y(_01317_));
 sky130_fd_sc_hd__nor2_2 _17211_ (.A(_11700_),
    .B(_12093_),
    .Y(_01319_));
 sky130_fd_sc_hd__nor2_2 _17212_ (.A(_11700_),
    .B(_12097_),
    .Y(_01321_));
 sky130_fd_sc_hd__nor2_2 _17213_ (.A(_11700_),
    .B(_12101_),
    .Y(_01323_));
 sky130_fd_sc_hd__buf_1 _17214_ (.A(is_slli_srli_srai),
    .X(_12432_));
 sky130_fd_sc_hd__buf_1 _17215_ (.A(_12432_),
    .X(_12433_));
 sky130_fd_sc_hd__nor2_2 _17216_ (.A(_12433_),
    .B(_12105_),
    .Y(_01325_));
 sky130_fd_sc_hd__nor2_2 _17217_ (.A(_12433_),
    .B(_12111_),
    .Y(_01327_));
 sky130_fd_sc_hd__nor2_2 _17218_ (.A(_12433_),
    .B(_12115_),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2_2 _17219_ (.A(_12433_),
    .B(_12122_),
    .Y(_01331_));
 sky130_fd_sc_hd__nor2_2 _17220_ (.A(_12433_),
    .B(_12126_),
    .Y(_01333_));
 sky130_fd_sc_hd__nor2_2 _17221_ (.A(_12433_),
    .B(_12129_),
    .Y(_01335_));
 sky130_fd_sc_hd__buf_1 _17222_ (.A(_12432_),
    .X(_12434_));
 sky130_fd_sc_hd__nor2_2 _17223_ (.A(_12434_),
    .B(_12134_),
    .Y(_01337_));
 sky130_fd_sc_hd__nor2_2 _17224_ (.A(_12434_),
    .B(_12138_),
    .Y(_01339_));
 sky130_fd_sc_hd__nor2_2 _17225_ (.A(_12434_),
    .B(_12142_),
    .Y(_01341_));
 sky130_fd_sc_hd__nor2_2 _17226_ (.A(_12434_),
    .B(_12146_),
    .Y(_01343_));
 sky130_vsdinv _17227_ (.A(\decoded_imm[20] ),
    .Y(_12435_));
 sky130_fd_sc_hd__nor2_2 _17228_ (.A(_12434_),
    .B(_12435_),
    .Y(_01345_));
 sky130_vsdinv _17229_ (.A(\decoded_imm[21] ),
    .Y(_12436_));
 sky130_fd_sc_hd__nor2_2 _17230_ (.A(_12434_),
    .B(_12436_),
    .Y(_01347_));
 sky130_fd_sc_hd__buf_1 _17231_ (.A(is_slli_srli_srai),
    .X(_12437_));
 sky130_vsdinv _17232_ (.A(\decoded_imm[22] ),
    .Y(_12438_));
 sky130_fd_sc_hd__nor2_2 _17233_ (.A(_12437_),
    .B(_12438_),
    .Y(_01349_));
 sky130_vsdinv _17234_ (.A(\decoded_imm[23] ),
    .Y(_12439_));
 sky130_fd_sc_hd__nor2_2 _17235_ (.A(_12437_),
    .B(_12439_),
    .Y(_01351_));
 sky130_vsdinv _17236_ (.A(\decoded_imm[24] ),
    .Y(_12440_));
 sky130_fd_sc_hd__nor2_2 _17237_ (.A(_12437_),
    .B(_12440_),
    .Y(_01353_));
 sky130_vsdinv _17238_ (.A(\decoded_imm[25] ),
    .Y(_12441_));
 sky130_fd_sc_hd__nor2_2 _17239_ (.A(_12437_),
    .B(_12441_),
    .Y(_01355_));
 sky130_vsdinv _17240_ (.A(\decoded_imm[26] ),
    .Y(_12442_));
 sky130_fd_sc_hd__nor2_2 _17241_ (.A(_12437_),
    .B(_12442_),
    .Y(_01357_));
 sky130_vsdinv _17242_ (.A(\decoded_imm[27] ),
    .Y(_12443_));
 sky130_fd_sc_hd__nor2_2 _17243_ (.A(_12437_),
    .B(_12443_),
    .Y(_01359_));
 sky130_vsdinv _17244_ (.A(\decoded_imm[28] ),
    .Y(_12444_));
 sky130_fd_sc_hd__nor2_2 _17245_ (.A(_12432_),
    .B(_12444_),
    .Y(_01361_));
 sky130_vsdinv _17246_ (.A(\decoded_imm[29] ),
    .Y(_12445_));
 sky130_fd_sc_hd__nor2_2 _17247_ (.A(_12432_),
    .B(_12445_),
    .Y(_01363_));
 sky130_vsdinv _17248_ (.A(\decoded_imm[30] ),
    .Y(_12446_));
 sky130_fd_sc_hd__nor2_2 _17249_ (.A(_12432_),
    .B(_12446_),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2_2 _17250_ (.A(_12432_),
    .B(_12173_),
    .Y(_01367_));
 sky130_vsdinv _17251_ (.A(\reg_next_pc[0] ),
    .Y(_12447_));
 sky130_fd_sc_hd__nor2_2 _17252_ (.A(_11797_),
    .B(_12447_),
    .Y(_01369_));
 sky130_fd_sc_hd__nor2_2 _17253_ (.A(_11715_),
    .B(_12195_),
    .Y(_12448_));
 sky130_fd_sc_hd__a21oi_2 _17254_ (.A1(_11715_),
    .A2(_12196_),
    .B1(_12448_),
    .Y(_01371_));
 sky130_vsdinv _17255_ (.A(\reg_pc[1] ),
    .Y(_12449_));
 sky130_fd_sc_hd__buf_1 _17256_ (.A(_11797_),
    .X(_12450_));
 sky130_fd_sc_hd__nor2_2 _17257_ (.A(_12449_),
    .B(_12450_),
    .Y(_01372_));
 sky130_vsdinv _17258_ (.A(pcpi_rs1[1]),
    .Y(_12451_));
 sky130_fd_sc_hd__o22a_2 _17259_ (.A1(_12451_),
    .A2(_12058_),
    .B1(_11861_),
    .B2(\decoded_imm[1] ),
    .X(_12452_));
 sky130_fd_sc_hd__o2bb2a_2 _17260_ (.A1_N(_12448_),
    .A2_N(_12452_),
    .B1(_12448_),
    .B2(_12452_),
    .X(_01374_));
 sky130_fd_sc_hd__inv_2 _17261_ (.A(\reg_pc[2] ),
    .Y(_02073_));
 sky130_fd_sc_hd__nor2_2 _17262_ (.A(_02073_),
    .B(_12450_),
    .Y(_01375_));
 sky130_fd_sc_hd__a22o_2 _17263_ (.A1(_11861_),
    .A2(\decoded_imm[1] ),
    .B1(_12448_),
    .B2(_12452_),
    .X(_12453_));
 sky130_fd_sc_hd__nor2_2 _17264_ (.A(pcpi_rs1[2]),
    .B(\decoded_imm[2] ),
    .Y(_12454_));
 sky130_fd_sc_hd__a21oi_2 _17265_ (.A1(_11860_),
    .A2(\decoded_imm[2] ),
    .B1(_12454_),
    .Y(_12455_));
 sky130_vsdinv _17266_ (.A(_12453_),
    .Y(_12456_));
 sky130_vsdinv _17267_ (.A(_12455_),
    .Y(_12457_));
 sky130_fd_sc_hd__o22a_2 _17268_ (.A1(_12453_),
    .A2(_12455_),
    .B1(_12456_),
    .B2(_12457_),
    .X(_01377_));
 sky130_vsdinv _17269_ (.A(\reg_pc[3] ),
    .Y(_12458_));
 sky130_fd_sc_hd__nor2_2 _17270_ (.A(_12458_),
    .B(_12450_),
    .Y(_01378_));
 sky130_vsdinv _17271_ (.A(pcpi_rs1[2]),
    .Y(_12459_));
 sky130_fd_sc_hd__o22a_2 _17272_ (.A1(_12459_),
    .A2(_12065_),
    .B1(_12456_),
    .B2(_12454_),
    .X(_12460_));
 sky130_fd_sc_hd__nor2_2 _17273_ (.A(pcpi_rs1[3]),
    .B(\decoded_imm[3] ),
    .Y(_12461_));
 sky130_fd_sc_hd__a21o_2 _17274_ (.A1(_11859_),
    .A2(\decoded_imm[3] ),
    .B1(_12461_),
    .X(_12462_));
 sky130_fd_sc_hd__o2bb2a_2 _17275_ (.A1_N(_12460_),
    .A2_N(_12462_),
    .B1(_12460_),
    .B2(_12462_),
    .X(_01380_));
 sky130_vsdinv _17276_ (.A(\reg_pc[4] ),
    .Y(_12463_));
 sky130_fd_sc_hd__nor2_2 _17277_ (.A(_12463_),
    .B(_12450_),
    .Y(_01381_));
 sky130_vsdinv _17278_ (.A(pcpi_rs1[3]),
    .Y(_12464_));
 sky130_fd_sc_hd__o22a_2 _17279_ (.A1(_12464_),
    .A2(_12071_),
    .B1(_12460_),
    .B2(_12461_),
    .X(_12465_));
 sky130_fd_sc_hd__nor2_2 _17280_ (.A(pcpi_rs1[4]),
    .B(\decoded_imm[4] ),
    .Y(_12466_));
 sky130_fd_sc_hd__a21o_2 _17281_ (.A1(_11858_),
    .A2(\decoded_imm[4] ),
    .B1(_12466_),
    .X(_12467_));
 sky130_fd_sc_hd__o2bb2a_2 _17282_ (.A1_N(_12465_),
    .A2_N(_12467_),
    .B1(_12465_),
    .B2(_12467_),
    .X(_01383_));
 sky130_vsdinv _17283_ (.A(\reg_pc[5] ),
    .Y(_12468_));
 sky130_fd_sc_hd__nor2_2 _17284_ (.A(_12468_),
    .B(_12450_),
    .Y(_01384_));
 sky130_vsdinv _17285_ (.A(pcpi_rs1[4]),
    .Y(_12469_));
 sky130_fd_sc_hd__o22a_2 _17286_ (.A1(_12469_),
    .A2(_12077_),
    .B1(_12465_),
    .B2(_12466_),
    .X(_12470_));
 sky130_fd_sc_hd__nor2_2 _17287_ (.A(pcpi_rs1[5]),
    .B(\decoded_imm[5] ),
    .Y(_12471_));
 sky130_fd_sc_hd__a21o_2 _17288_ (.A1(_11857_),
    .A2(\decoded_imm[5] ),
    .B1(_12471_),
    .X(_12472_));
 sky130_fd_sc_hd__o2bb2a_2 _17289_ (.A1_N(_12470_),
    .A2_N(_12472_),
    .B1(_12470_),
    .B2(_12472_),
    .X(_01386_));
 sky130_vsdinv _17290_ (.A(\reg_pc[6] ),
    .Y(_12473_));
 sky130_fd_sc_hd__nor2_2 _17291_ (.A(_12473_),
    .B(_12450_),
    .Y(_01387_));
 sky130_vsdinv _17292_ (.A(pcpi_rs1[5]),
    .Y(_12474_));
 sky130_fd_sc_hd__o22ai_2 _17293_ (.A1(_12474_),
    .A2(_12084_),
    .B1(_12470_),
    .B2(_12471_),
    .Y(_12475_));
 sky130_vsdinv _17294_ (.A(pcpi_rs1[6]),
    .Y(_12476_));
 sky130_fd_sc_hd__o22a_2 _17295_ (.A1(_12476_),
    .A2(_12091_),
    .B1(_11855_),
    .B2(\decoded_imm[6] ),
    .X(_12477_));
 sky130_fd_sc_hd__o2bb2a_2 _17296_ (.A1_N(_12475_),
    .A2_N(_12477_),
    .B1(_12475_),
    .B2(_12477_),
    .X(_01389_));
 sky130_vsdinv _17297_ (.A(\reg_pc[7] ),
    .Y(_12478_));
 sky130_fd_sc_hd__buf_1 _17298_ (.A(_11797_),
    .X(_12479_));
 sky130_fd_sc_hd__nor2_2 _17299_ (.A(_12478_),
    .B(_12479_),
    .Y(_01390_));
 sky130_fd_sc_hd__nor2_2 _17300_ (.A(pcpi_rs1[7]),
    .B(\decoded_imm[7] ),
    .Y(_12480_));
 sky130_fd_sc_hd__a21oi_2 _17301_ (.A1(_11852_),
    .A2(\decoded_imm[7] ),
    .B1(_12480_),
    .Y(_12481_));
 sky130_fd_sc_hd__a22o_2 _17302_ (.A1(_11856_),
    .A2(\decoded_imm[6] ),
    .B1(_12475_),
    .B2(_12477_),
    .X(_12482_));
 sky130_fd_sc_hd__a2bb2oi_2 _17303_ (.A1_N(_12481_),
    .A2_N(_12482_),
    .B1(_12481_),
    .B2(_12482_),
    .Y(_01392_));
 sky130_vsdinv _17304_ (.A(\reg_pc[8] ),
    .Y(_12483_));
 sky130_fd_sc_hd__nor2_2 _17305_ (.A(_12483_),
    .B(_12479_),
    .Y(_01393_));
 sky130_vsdinv _17306_ (.A(_11852_),
    .Y(_12484_));
 sky130_fd_sc_hd__o32a_2 _17307_ (.A1(_12476_),
    .A2(_12091_),
    .A3(_12480_),
    .B1(_12484_),
    .B2(_12093_),
    .X(_12485_));
 sky130_vsdinv _17308_ (.A(_12485_),
    .Y(_12486_));
 sky130_fd_sc_hd__a31o_2 _17309_ (.A1(_12477_),
    .A2(_12481_),
    .A3(_12475_),
    .B1(_12486_),
    .X(_12487_));
 sky130_vsdinv _17310_ (.A(_12487_),
    .Y(_12488_));
 sky130_vsdinv _17311_ (.A(pcpi_rs1[8]),
    .Y(_12489_));
 sky130_fd_sc_hd__o22a_2 _17312_ (.A1(_12489_),
    .A2(_12097_),
    .B1(pcpi_rs1[8]),
    .B2(\decoded_imm[8] ),
    .X(_12490_));
 sky130_vsdinv _17313_ (.A(_12490_),
    .Y(_12491_));
 sky130_fd_sc_hd__o22a_2 _17314_ (.A1(_12488_),
    .A2(_12491_),
    .B1(_12487_),
    .B2(_12490_),
    .X(_01395_));
 sky130_vsdinv _17315_ (.A(\reg_pc[9] ),
    .Y(_12492_));
 sky130_fd_sc_hd__nor2_2 _17316_ (.A(_12492_),
    .B(_12479_),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_2 _17317_ (.A(_11848_),
    .B(\decoded_imm[9] ),
    .Y(_12493_));
 sky130_fd_sc_hd__a21o_2 _17318_ (.A1(_11848_),
    .A2(\decoded_imm[9] ),
    .B1(_12493_),
    .X(_12494_));
 sky130_fd_sc_hd__o22a_2 _17319_ (.A1(_12489_),
    .A2(_12097_),
    .B1(_12488_),
    .B2(_12491_),
    .X(_12495_));
 sky130_fd_sc_hd__o2bb2a_2 _17320_ (.A1_N(_12494_),
    .A2_N(_12495_),
    .B1(_12494_),
    .B2(_12495_),
    .X(_01398_));
 sky130_vsdinv _17321_ (.A(\reg_pc[10] ),
    .Y(_12496_));
 sky130_fd_sc_hd__nor2_2 _17322_ (.A(_12496_),
    .B(_12479_),
    .Y(_01399_));
 sky130_vsdinv _17323_ (.A(pcpi_rs1[10]),
    .Y(_12497_));
 sky130_fd_sc_hd__a22o_2 _17324_ (.A1(pcpi_rs1[10]),
    .A2(\decoded_imm[10] ),
    .B1(_12497_),
    .B2(_12105_),
    .X(_12498_));
 sky130_vsdinv _17325_ (.A(_11848_),
    .Y(_12499_));
 sky130_fd_sc_hd__o32a_2 _17326_ (.A1(_12489_),
    .A2(_12097_),
    .A3(_12493_),
    .B1(_12499_),
    .B2(_12101_),
    .X(_12500_));
 sky130_fd_sc_hd__o31a_2 _17327_ (.A1(_12491_),
    .A2(_12494_),
    .A3(_12488_),
    .B1(_12500_),
    .X(_12501_));
 sky130_fd_sc_hd__a2bb2oi_2 _17328_ (.A1_N(_12498_),
    .A2_N(_12501_),
    .B1(_12498_),
    .B2(_12501_),
    .Y(_01401_));
 sky130_vsdinv _17329_ (.A(\reg_pc[11] ),
    .Y(_12502_));
 sky130_fd_sc_hd__nor2_2 _17330_ (.A(_12502_),
    .B(_12479_),
    .Y(_01402_));
 sky130_vsdinv _17331_ (.A(pcpi_rs1[11]),
    .Y(_12503_));
 sky130_fd_sc_hd__a22o_2 _17332_ (.A1(pcpi_rs1[11]),
    .A2(\decoded_imm[11] ),
    .B1(_12503_),
    .B2(_12111_),
    .X(_12504_));
 sky130_fd_sc_hd__o22a_2 _17333_ (.A1(_12497_),
    .A2(_12105_),
    .B1(_12498_),
    .B2(_12501_),
    .X(_12505_));
 sky130_fd_sc_hd__a2bb2oi_2 _17334_ (.A1_N(_12504_),
    .A2_N(_12505_),
    .B1(_12504_),
    .B2(_12505_),
    .Y(_01404_));
 sky130_vsdinv _17335_ (.A(\reg_pc[12] ),
    .Y(_12506_));
 sky130_fd_sc_hd__nor2_2 _17336_ (.A(_12506_),
    .B(_12479_),
    .Y(_01405_));
 sky130_vsdinv _17337_ (.A(pcpi_rs1[12]),
    .Y(_12507_));
 sky130_fd_sc_hd__a22o_2 _17338_ (.A1(pcpi_rs1[12]),
    .A2(\decoded_imm[12] ),
    .B1(_12507_),
    .B2(_12115_),
    .X(_12508_));
 sky130_fd_sc_hd__o22a_2 _17339_ (.A1(_12503_),
    .A2(_12111_),
    .B1(_12504_),
    .B2(_12505_),
    .X(_12509_));
 sky130_fd_sc_hd__a2bb2oi_2 _17340_ (.A1_N(_12508_),
    .A2_N(_12509_),
    .B1(_12508_),
    .B2(_12509_),
    .Y(_01407_));
 sky130_vsdinv _17341_ (.A(\reg_pc[13] ),
    .Y(_12510_));
 sky130_fd_sc_hd__buf_1 _17342_ (.A(_11797_),
    .X(_12511_));
 sky130_fd_sc_hd__nor2_2 _17343_ (.A(_12510_),
    .B(_12511_),
    .Y(_01408_));
 sky130_vsdinv _17344_ (.A(pcpi_rs1[13]),
    .Y(_12512_));
 sky130_fd_sc_hd__a22o_2 _17345_ (.A1(pcpi_rs1[13]),
    .A2(\decoded_imm[13] ),
    .B1(_12512_),
    .B2(_12122_),
    .X(_12513_));
 sky130_fd_sc_hd__o22a_2 _17346_ (.A1(_12507_),
    .A2(_12115_),
    .B1(_12508_),
    .B2(_12509_),
    .X(_12514_));
 sky130_fd_sc_hd__a2bb2oi_2 _17347_ (.A1_N(_12513_),
    .A2_N(_12514_),
    .B1(_12513_),
    .B2(_12514_),
    .Y(_01410_));
 sky130_vsdinv _17348_ (.A(\reg_pc[14] ),
    .Y(_12515_));
 sky130_fd_sc_hd__nor2_2 _17349_ (.A(_12515_),
    .B(_12511_),
    .Y(_01411_));
 sky130_vsdinv _17350_ (.A(pcpi_rs1[14]),
    .Y(_12516_));
 sky130_fd_sc_hd__a22o_2 _17351_ (.A1(pcpi_rs1[14]),
    .A2(\decoded_imm[14] ),
    .B1(_12516_),
    .B2(_12126_),
    .X(_12517_));
 sky130_fd_sc_hd__o22a_2 _17352_ (.A1(_12512_),
    .A2(_12122_),
    .B1(_12513_),
    .B2(_12514_),
    .X(_12518_));
 sky130_fd_sc_hd__a2bb2oi_2 _17353_ (.A1_N(_12517_),
    .A2_N(_12518_),
    .B1(_12517_),
    .B2(_12518_),
    .Y(_01413_));
 sky130_vsdinv _17354_ (.A(\reg_pc[15] ),
    .Y(_12519_));
 sky130_fd_sc_hd__nor2_2 _17355_ (.A(_12519_),
    .B(_12511_),
    .Y(_01414_));
 sky130_vsdinv _17356_ (.A(pcpi_rs1[15]),
    .Y(_12520_));
 sky130_fd_sc_hd__a22o_2 _17357_ (.A1(pcpi_rs1[15]),
    .A2(\decoded_imm[15] ),
    .B1(_12520_),
    .B2(_12129_),
    .X(_12521_));
 sky130_fd_sc_hd__o22a_2 _17358_ (.A1(_12516_),
    .A2(_12126_),
    .B1(_12517_),
    .B2(_12518_),
    .X(_12522_));
 sky130_fd_sc_hd__a2bb2oi_2 _17359_ (.A1_N(_12521_),
    .A2_N(_12522_),
    .B1(_12521_),
    .B2(_12522_),
    .Y(_01416_));
 sky130_vsdinv _17360_ (.A(\reg_pc[16] ),
    .Y(_12523_));
 sky130_fd_sc_hd__nor2_2 _17361_ (.A(_12523_),
    .B(_12511_),
    .Y(_01417_));
 sky130_fd_sc_hd__o22a_2 _17362_ (.A1(_12520_),
    .A2(_12129_),
    .B1(_12521_),
    .B2(_12522_),
    .X(_12524_));
 sky130_vsdinv _17363_ (.A(pcpi_rs1[16]),
    .Y(_12525_));
 sky130_fd_sc_hd__o22a_2 _17364_ (.A1(_12525_),
    .A2(_12134_),
    .B1(pcpi_rs1[16]),
    .B2(\decoded_imm[16] ),
    .X(_12526_));
 sky130_vsdinv _17365_ (.A(_12526_),
    .Y(_12527_));
 sky130_vsdinv _17366_ (.A(_12524_),
    .Y(_12528_));
 sky130_fd_sc_hd__o22a_2 _17367_ (.A1(_12524_),
    .A2(_12527_),
    .B1(_12528_),
    .B2(_12526_),
    .X(_01419_));
 sky130_vsdinv _17368_ (.A(\reg_pc[17] ),
    .Y(_12529_));
 sky130_fd_sc_hd__nor2_2 _17369_ (.A(_12529_),
    .B(_12511_),
    .Y(_01420_));
 sky130_fd_sc_hd__nor2_2 _17370_ (.A(_11837_),
    .B(\decoded_imm[17] ),
    .Y(_12530_));
 sky130_fd_sc_hd__a21o_2 _17371_ (.A1(_11837_),
    .A2(\decoded_imm[17] ),
    .B1(_12530_),
    .X(_12531_));
 sky130_fd_sc_hd__o22a_2 _17372_ (.A1(_12525_),
    .A2(_12134_),
    .B1(_12524_),
    .B2(_12527_),
    .X(_12532_));
 sky130_fd_sc_hd__o2bb2a_2 _17373_ (.A1_N(_12531_),
    .A2_N(_12532_),
    .B1(_12531_),
    .B2(_12532_),
    .X(_01422_));
 sky130_vsdinv _17374_ (.A(\reg_pc[18] ),
    .Y(_12533_));
 sky130_fd_sc_hd__nor2_2 _17375_ (.A(_12533_),
    .B(_12511_),
    .Y(_01423_));
 sky130_vsdinv _17376_ (.A(pcpi_rs1[18]),
    .Y(_12534_));
 sky130_fd_sc_hd__a22o_2 _17377_ (.A1(_11836_),
    .A2(\decoded_imm[18] ),
    .B1(_12534_),
    .B2(_12142_),
    .X(_12535_));
 sky130_vsdinv _17378_ (.A(_11837_),
    .Y(_12536_));
 sky130_fd_sc_hd__o32a_2 _17379_ (.A1(_12525_),
    .A2(_12134_),
    .A3(_12530_),
    .B1(_12536_),
    .B2(_12138_),
    .X(_12537_));
 sky130_fd_sc_hd__o31a_2 _17380_ (.A1(_12527_),
    .A2(_12531_),
    .A3(_12524_),
    .B1(_12537_),
    .X(_12538_));
 sky130_fd_sc_hd__a2bb2oi_2 _17381_ (.A1_N(_12535_),
    .A2_N(_12538_),
    .B1(_12535_),
    .B2(_12538_),
    .Y(_01425_));
 sky130_vsdinv _17382_ (.A(\reg_pc[19] ),
    .Y(_12539_));
 sky130_fd_sc_hd__buf_1 _17383_ (.A(instr_lui),
    .X(_12540_));
 sky130_fd_sc_hd__nor2_2 _17384_ (.A(_12539_),
    .B(_12540_),
    .Y(_01426_));
 sky130_vsdinv _17385_ (.A(pcpi_rs1[19]),
    .Y(_12541_));
 sky130_fd_sc_hd__a22o_2 _17386_ (.A1(_11834_),
    .A2(\decoded_imm[19] ),
    .B1(_12541_),
    .B2(_12146_),
    .X(_12542_));
 sky130_fd_sc_hd__o22a_2 _17387_ (.A1(_12534_),
    .A2(_12142_),
    .B1(_12535_),
    .B2(_12538_),
    .X(_12543_));
 sky130_fd_sc_hd__a2bb2oi_2 _17388_ (.A1_N(_12542_),
    .A2_N(_12543_),
    .B1(_12542_),
    .B2(_12543_),
    .Y(_01428_));
 sky130_vsdinv _17389_ (.A(\reg_pc[20] ),
    .Y(_12544_));
 sky130_fd_sc_hd__nor2_2 _17390_ (.A(_12544_),
    .B(_12540_),
    .Y(_01429_));
 sky130_vsdinv _17391_ (.A(pcpi_rs1[20]),
    .Y(_12545_));
 sky130_fd_sc_hd__a22o_2 _17392_ (.A1(_11832_),
    .A2(\decoded_imm[20] ),
    .B1(_12545_),
    .B2(_12435_),
    .X(_12546_));
 sky130_fd_sc_hd__o22a_2 _17393_ (.A1(_12541_),
    .A2(_12146_),
    .B1(_12542_),
    .B2(_12543_),
    .X(_12547_));
 sky130_fd_sc_hd__a2bb2oi_2 _17394_ (.A1_N(_12546_),
    .A2_N(_12547_),
    .B1(_12546_),
    .B2(_12547_),
    .Y(_01431_));
 sky130_vsdinv _17395_ (.A(\reg_pc[21] ),
    .Y(_12548_));
 sky130_fd_sc_hd__nor2_2 _17396_ (.A(_12548_),
    .B(_12540_),
    .Y(_01432_));
 sky130_vsdinv _17397_ (.A(pcpi_rs1[21]),
    .Y(_12549_));
 sky130_fd_sc_hd__a22o_2 _17398_ (.A1(_11831_),
    .A2(\decoded_imm[21] ),
    .B1(_12549_),
    .B2(_12436_),
    .X(_12550_));
 sky130_fd_sc_hd__o22a_2 _17399_ (.A1(_12545_),
    .A2(_12435_),
    .B1(_12546_),
    .B2(_12547_),
    .X(_12551_));
 sky130_fd_sc_hd__a2bb2oi_2 _17400_ (.A1_N(_12550_),
    .A2_N(_12551_),
    .B1(_12550_),
    .B2(_12551_),
    .Y(_01434_));
 sky130_vsdinv _17401_ (.A(\reg_pc[22] ),
    .Y(_12552_));
 sky130_fd_sc_hd__nor2_2 _17402_ (.A(_12552_),
    .B(_12540_),
    .Y(_01435_));
 sky130_vsdinv _17403_ (.A(pcpi_rs1[22]),
    .Y(_12553_));
 sky130_fd_sc_hd__a22o_2 _17404_ (.A1(_11830_),
    .A2(\decoded_imm[22] ),
    .B1(_12553_),
    .B2(_12438_),
    .X(_12554_));
 sky130_fd_sc_hd__o22a_2 _17405_ (.A1(_12549_),
    .A2(_12436_),
    .B1(_12550_),
    .B2(_12551_),
    .X(_12555_));
 sky130_fd_sc_hd__a2bb2oi_2 _17406_ (.A1_N(_12554_),
    .A2_N(_12555_),
    .B1(_12554_),
    .B2(_12555_),
    .Y(_01437_));
 sky130_vsdinv _17407_ (.A(\reg_pc[23] ),
    .Y(_12556_));
 sky130_fd_sc_hd__nor2_2 _17408_ (.A(_12556_),
    .B(_12540_),
    .Y(_01438_));
 sky130_vsdinv _17409_ (.A(pcpi_rs1[23]),
    .Y(_12557_));
 sky130_fd_sc_hd__a22o_2 _17410_ (.A1(_11829_),
    .A2(\decoded_imm[23] ),
    .B1(_12557_),
    .B2(_12439_),
    .X(_12558_));
 sky130_fd_sc_hd__o22a_2 _17411_ (.A1(_12553_),
    .A2(_12438_),
    .B1(_12554_),
    .B2(_12555_),
    .X(_12559_));
 sky130_fd_sc_hd__a2bb2oi_2 _17412_ (.A1_N(_12558_),
    .A2_N(_12559_),
    .B1(_12558_),
    .B2(_12559_),
    .Y(_01440_));
 sky130_vsdinv _17413_ (.A(\reg_pc[24] ),
    .Y(_12560_));
 sky130_fd_sc_hd__nor2_2 _17414_ (.A(_12560_),
    .B(_12540_),
    .Y(_01441_));
 sky130_fd_sc_hd__o22ai_2 _17415_ (.A1(_12557_),
    .A2(_12439_),
    .B1(_12558_),
    .B2(_12559_),
    .Y(_12561_));
 sky130_vsdinv _17416_ (.A(_11827_),
    .Y(_12562_));
 sky130_fd_sc_hd__o22a_2 _17417_ (.A1(_12562_),
    .A2(_12440_),
    .B1(_11827_),
    .B2(\decoded_imm[24] ),
    .X(_12563_));
 sky130_fd_sc_hd__o2bb2a_2 _17418_ (.A1_N(_12561_),
    .A2_N(_12563_),
    .B1(_12561_),
    .B2(_12563_),
    .X(_01443_));
 sky130_vsdinv _17419_ (.A(\reg_pc[25] ),
    .Y(_12564_));
 sky130_fd_sc_hd__buf_1 _17420_ (.A(instr_lui),
    .X(_12565_));
 sky130_fd_sc_hd__nor2_2 _17421_ (.A(_12564_),
    .B(_12565_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_2 _17422_ (.A(_11824_),
    .B(\decoded_imm[25] ),
    .Y(_12566_));
 sky130_fd_sc_hd__a21oi_2 _17423_ (.A1(_11825_),
    .A2(\decoded_imm[25] ),
    .B1(_12566_),
    .Y(_12567_));
 sky130_fd_sc_hd__a22o_2 _17424_ (.A1(_11828_),
    .A2(\decoded_imm[24] ),
    .B1(_12561_),
    .B2(_12563_),
    .X(_12568_));
 sky130_fd_sc_hd__a2bb2oi_2 _17425_ (.A1_N(_12567_),
    .A2_N(_12568_),
    .B1(_12567_),
    .B2(_12568_),
    .Y(_01446_));
 sky130_vsdinv _17426_ (.A(\reg_pc[26] ),
    .Y(_12569_));
 sky130_fd_sc_hd__nor2_2 _17427_ (.A(_12569_),
    .B(_12565_),
    .Y(_01447_));
 sky130_vsdinv _17428_ (.A(_11824_),
    .Y(_12570_));
 sky130_fd_sc_hd__o32a_2 _17429_ (.A1(_12562_),
    .A2(_12440_),
    .A3(_12566_),
    .B1(_12570_),
    .B2(_12441_),
    .X(_12571_));
 sky130_vsdinv _17430_ (.A(_12571_),
    .Y(_12572_));
 sky130_fd_sc_hd__a31o_2 _17431_ (.A1(_12563_),
    .A2(_12567_),
    .A3(_12561_),
    .B1(_12572_),
    .X(_12573_));
 sky130_vsdinv _17432_ (.A(_11821_),
    .Y(_12574_));
 sky130_fd_sc_hd__o22a_2 _17433_ (.A1(_12574_),
    .A2(_12442_),
    .B1(_11822_),
    .B2(\decoded_imm[26] ),
    .X(_12575_));
 sky130_fd_sc_hd__o2bb2a_2 _17434_ (.A1_N(_12573_),
    .A2_N(_12575_),
    .B1(_12573_),
    .B2(_12575_),
    .X(_01449_));
 sky130_vsdinv _17435_ (.A(\reg_pc[27] ),
    .Y(_12576_));
 sky130_fd_sc_hd__nor2_2 _17436_ (.A(_12576_),
    .B(_12565_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_2 _17437_ (.A(_11819_),
    .B(\decoded_imm[27] ),
    .Y(_12577_));
 sky130_fd_sc_hd__a21oi_2 _17438_ (.A1(_11820_),
    .A2(\decoded_imm[27] ),
    .B1(_12577_),
    .Y(_12578_));
 sky130_fd_sc_hd__a22o_2 _17439_ (.A1(_11822_),
    .A2(\decoded_imm[26] ),
    .B1(_12573_),
    .B2(_12575_),
    .X(_12579_));
 sky130_fd_sc_hd__a2bb2oi_2 _17440_ (.A1_N(_12578_),
    .A2_N(_12579_),
    .B1(_12578_),
    .B2(_12579_),
    .Y(_01452_));
 sky130_vsdinv _17441_ (.A(\reg_pc[28] ),
    .Y(_12580_));
 sky130_fd_sc_hd__nor2_2 _17442_ (.A(_12580_),
    .B(_12565_),
    .Y(_01453_));
 sky130_vsdinv _17443_ (.A(_11819_),
    .Y(_12581_));
 sky130_fd_sc_hd__o32a_2 _17444_ (.A1(_12574_),
    .A2(_12442_),
    .A3(_12577_),
    .B1(_12581_),
    .B2(_12443_),
    .X(_12582_));
 sky130_vsdinv _17445_ (.A(_12582_),
    .Y(_12583_));
 sky130_fd_sc_hd__a31o_2 _17446_ (.A1(_12575_),
    .A2(_12578_),
    .A3(_12573_),
    .B1(_12583_),
    .X(_12584_));
 sky130_fd_sc_hd__nor2_2 _17447_ (.A(pcpi_rs1[28]),
    .B(\decoded_imm[28] ),
    .Y(_12585_));
 sky130_fd_sc_hd__a21oi_2 _17448_ (.A1(_11818_),
    .A2(\decoded_imm[28] ),
    .B1(_12585_),
    .Y(_12586_));
 sky130_vsdinv _17449_ (.A(_12584_),
    .Y(_12587_));
 sky130_vsdinv _17450_ (.A(_12586_),
    .Y(_12588_));
 sky130_fd_sc_hd__o22a_2 _17451_ (.A1(_12584_),
    .A2(_12586_),
    .B1(_12587_),
    .B2(_12588_),
    .X(_01455_));
 sky130_vsdinv _17452_ (.A(\reg_pc[29] ),
    .Y(_12589_));
 sky130_fd_sc_hd__nor2_2 _17453_ (.A(_12589_),
    .B(_12565_),
    .Y(_01456_));
 sky130_vsdinv _17454_ (.A(_11818_),
    .Y(_12590_));
 sky130_fd_sc_hd__o22a_2 _17455_ (.A1(_12590_),
    .A2(_12444_),
    .B1(_12587_),
    .B2(_12585_),
    .X(_12591_));
 sky130_fd_sc_hd__nor2_2 _17456_ (.A(_11817_),
    .B(\decoded_imm[29] ),
    .Y(_12592_));
 sky130_fd_sc_hd__a21o_2 _17457_ (.A1(_11817_),
    .A2(\decoded_imm[29] ),
    .B1(_12592_),
    .X(_12593_));
 sky130_fd_sc_hd__o2bb2a_2 _17458_ (.A1_N(_12591_),
    .A2_N(_12593_),
    .B1(_12591_),
    .B2(_12593_),
    .X(_01458_));
 sky130_vsdinv _17459_ (.A(\reg_pc[30] ),
    .Y(_12594_));
 sky130_fd_sc_hd__nor2_2 _17460_ (.A(_12594_),
    .B(_12565_),
    .Y(_01459_));
 sky130_vsdinv _17461_ (.A(_11816_),
    .Y(_12595_));
 sky130_fd_sc_hd__a22o_2 _17462_ (.A1(_11816_),
    .A2(\decoded_imm[30] ),
    .B1(_12595_),
    .B2(_12446_),
    .X(_12596_));
 sky130_vsdinv _17463_ (.A(pcpi_rs1[29]),
    .Y(_12597_));
 sky130_fd_sc_hd__o22a_2 _17464_ (.A1(_12597_),
    .A2(_12445_),
    .B1(_12591_),
    .B2(_12592_),
    .X(_12598_));
 sky130_fd_sc_hd__a2bb2oi_2 _17465_ (.A1_N(_12596_),
    .A2_N(_12598_),
    .B1(_12596_),
    .B2(_12598_),
    .Y(_01461_));
 sky130_vsdinv _17466_ (.A(\reg_pc[31] ),
    .Y(_12599_));
 sky130_fd_sc_hd__nor2_2 _17467_ (.A(_12599_),
    .B(_11797_),
    .Y(_01462_));
 sky130_fd_sc_hd__o22a_2 _17468_ (.A1(_12595_),
    .A2(_12446_),
    .B1(_12596_),
    .B2(_12598_),
    .X(_12600_));
 sky130_fd_sc_hd__o22a_2 _17469_ (.A1(_11812_),
    .A2(\decoded_imm[31] ),
    .B1(_10568_),
    .B2(_12173_),
    .X(_12601_));
 sky130_fd_sc_hd__o2bb2ai_2 _17470_ (.A1_N(_12600_),
    .A2_N(_12601_),
    .B1(_12600_),
    .B2(_12601_),
    .Y(_01464_));
 sky130_fd_sc_hd__and2_2 _17471_ (.A(_12376_),
    .B(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__and2_2 _17472_ (.A(_12376_),
    .B(_01469_),
    .X(_01470_));
 sky130_vsdinv _17473_ (.A(\reg_next_pc[4] ),
    .Y(_01471_));
 sky130_fd_sc_hd__a21oi_2 _17474_ (.A1(_12376_),
    .A2(_01473_),
    .B1(_10656_),
    .Y(_01474_));
 sky130_fd_sc_hd__and2_2 _17475_ (.A(_12376_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__and2_2 _17476_ (.A(_12376_),
    .B(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__buf_1 _17477_ (.A(_10473_),
    .X(_12602_));
 sky130_fd_sc_hd__and2_2 _17478_ (.A(_12602_),
    .B(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__and2_2 _17479_ (.A(_12602_),
    .B(_01486_),
    .X(_01487_));
 sky130_fd_sc_hd__and2_2 _17480_ (.A(_12602_),
    .B(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__and2_2 _17481_ (.A(_12602_),
    .B(_01492_),
    .X(_01493_));
 sky130_fd_sc_hd__and2_2 _17482_ (.A(_12602_),
    .B(_01495_),
    .X(_01496_));
 sky130_fd_sc_hd__and2_2 _17483_ (.A(_12602_),
    .B(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__buf_1 _17484_ (.A(_10473_),
    .X(_12603_));
 sky130_fd_sc_hd__and2_2 _17485_ (.A(_12603_),
    .B(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__and2_2 _17486_ (.A(_12603_),
    .B(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__and2_2 _17487_ (.A(_12603_),
    .B(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__and2_2 _17488_ (.A(_12603_),
    .B(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__and2_2 _17489_ (.A(_12603_),
    .B(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__and2_2 _17490_ (.A(_12603_),
    .B(_01516_),
    .X(_01517_));
 sky130_fd_sc_hd__buf_1 _17491_ (.A(_10473_),
    .X(_12604_));
 sky130_fd_sc_hd__and2_2 _17492_ (.A(_12604_),
    .B(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__and2_2 _17493_ (.A(_12604_),
    .B(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__and2_2 _17494_ (.A(_12604_),
    .B(_01525_),
    .X(_01526_));
 sky130_fd_sc_hd__and2_2 _17495_ (.A(_12604_),
    .B(_01528_),
    .X(_01529_));
 sky130_fd_sc_hd__and2_2 _17496_ (.A(_12604_),
    .B(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__and2_2 _17497_ (.A(_12604_),
    .B(_01534_),
    .X(_01535_));
 sky130_fd_sc_hd__buf_1 _17498_ (.A(latched_branch),
    .X(_12605_));
 sky130_fd_sc_hd__and2_2 _17499_ (.A(_12605_),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__and2_2 _17500_ (.A(_12605_),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__and2_2 _17501_ (.A(_12605_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__and2_2 _17502_ (.A(_12605_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__and2_2 _17503_ (.A(_12605_),
    .B(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__and2_2 _17504_ (.A(_12605_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__and2_2 _17505_ (.A(_10473_),
    .B(_01555_),
    .X(_01556_));
 sky130_vsdinv _17506_ (.A(_02590_),
    .Y(_12606_));
 sky130_fd_sc_hd__nor2_2 _17507_ (.A(_12606_),
    .B(_12061_),
    .Y(_12607_));
 sky130_fd_sc_hd__a21oi_2 _17508_ (.A1(_12606_),
    .A2(_12061_),
    .B1(_12607_),
    .Y(_01557_));
 sky130_fd_sc_hd__inv_2 _17509_ (.A(_02560_),
    .Y(_01561_));
 sky130_fd_sc_hd__o22a_2 _17510_ (.A1(_01561_),
    .A2(_12068_),
    .B1(_02560_),
    .B2(\decoded_imm_uj[2] ),
    .X(_12608_));
 sky130_fd_sc_hd__o2bb2a_2 _17511_ (.A1_N(_12607_),
    .A2_N(_12608_),
    .B1(_12607_),
    .B2(_12608_),
    .X(_01562_));
 sky130_fd_sc_hd__o22a_2 _17512_ (.A1(_01561_),
    .A2(_02410_),
    .B1(_02560_),
    .B2(_11102_),
    .X(_01565_));
 sky130_vsdinv _17513_ (.A(_02571_),
    .Y(_12609_));
 sky130_fd_sc_hd__nor2_2 _17514_ (.A(_12609_),
    .B(_01561_),
    .Y(_12610_));
 sky130_fd_sc_hd__a21oi_2 _17515_ (.A1(_12609_),
    .A2(_01561_),
    .B1(_12610_),
    .Y(_01567_));
 sky130_fd_sc_hd__a22o_2 _17516_ (.A1(_02560_),
    .A2(\decoded_imm_uj[2] ),
    .B1(_12607_),
    .B2(_12608_),
    .X(_12611_));
 sky130_fd_sc_hd__nor2_2 _17517_ (.A(_02571_),
    .B(\decoded_imm_uj[3] ),
    .Y(_12612_));
 sky130_fd_sc_hd__a21oi_2 _17518_ (.A1(_02571_),
    .A2(\decoded_imm_uj[3] ),
    .B1(_12612_),
    .Y(_12613_));
 sky130_vsdinv _17519_ (.A(_12611_),
    .Y(_12614_));
 sky130_vsdinv _17520_ (.A(_12613_),
    .Y(_12615_));
 sky130_fd_sc_hd__o22a_2 _17521_ (.A1(_12611_),
    .A2(_12613_),
    .B1(_12614_),
    .B2(_12615_),
    .X(_01568_));
 sky130_fd_sc_hd__nand2_2 _17522_ (.A(_02582_),
    .B(_12610_),
    .Y(_12616_));
 sky130_fd_sc_hd__o21a_2 _17523_ (.A1(_02582_),
    .A2(_12610_),
    .B1(_12616_),
    .X(_01571_));
 sky130_fd_sc_hd__o22a_2 _17524_ (.A1(_12609_),
    .A2(_12074_),
    .B1(_12614_),
    .B2(_12612_),
    .X(_12617_));
 sky130_vsdinv _17525_ (.A(_12617_),
    .Y(_12618_));
 sky130_fd_sc_hd__nor2_2 _17526_ (.A(\decoded_imm_uj[4] ),
    .B(_02582_),
    .Y(_12619_));
 sky130_fd_sc_hd__a21o_2 _17527_ (.A1(\decoded_imm_uj[4] ),
    .A2(_02582_),
    .B1(_12619_),
    .X(_12620_));
 sky130_fd_sc_hd__a2bb2o_2 _17528_ (.A1_N(_12618_),
    .A2_N(_12620_),
    .B1(_12618_),
    .B2(_12620_),
    .X(_01572_));
 sky130_vsdinv _17529_ (.A(_02583_),
    .Y(_12621_));
 sky130_fd_sc_hd__nor2_2 _17530_ (.A(_12621_),
    .B(_12616_),
    .Y(_12622_));
 sky130_fd_sc_hd__a21oi_2 _17531_ (.A1(_12621_),
    .A2(_12616_),
    .B1(_12622_),
    .Y(_01575_));
 sky130_fd_sc_hd__o22a_2 _17532_ (.A1(_00367_),
    .A2(_01475_),
    .B1(_12617_),
    .B2(_12619_),
    .X(_12623_));
 sky130_fd_sc_hd__nor2_2 _17533_ (.A(_02583_),
    .B(\decoded_imm_uj[5] ),
    .Y(_12624_));
 sky130_fd_sc_hd__a21o_2 _17534_ (.A1(_02583_),
    .A2(\decoded_imm_uj[5] ),
    .B1(_12624_),
    .X(_12625_));
 sky130_fd_sc_hd__o2bb2a_2 _17535_ (.A1_N(_12623_),
    .A2_N(_12625_),
    .B1(_12623_),
    .B2(_12625_),
    .X(_01576_));
 sky130_fd_sc_hd__nand2_2 _17536_ (.A(_02584_),
    .B(_12622_),
    .Y(_12626_));
 sky130_fd_sc_hd__o21a_2 _17537_ (.A1(_02584_),
    .A2(_12622_),
    .B1(_12626_),
    .X(_01579_));
 sky130_fd_sc_hd__o22a_2 _17538_ (.A1(_12621_),
    .A2(_12085_),
    .B1(_12623_),
    .B2(_12624_),
    .X(_12627_));
 sky130_fd_sc_hd__nor2_2 _17539_ (.A(_02584_),
    .B(\decoded_imm_uj[6] ),
    .Y(_12628_));
 sky130_fd_sc_hd__a21o_2 _17540_ (.A1(_02584_),
    .A2(\decoded_imm_uj[6] ),
    .B1(_12628_),
    .X(_12629_));
 sky130_fd_sc_hd__o2bb2a_2 _17541_ (.A1_N(_12627_),
    .A2_N(_12629_),
    .B1(_12627_),
    .B2(_12629_),
    .X(_01580_));
 sky130_vsdinv _17542_ (.A(_02585_),
    .Y(_12630_));
 sky130_fd_sc_hd__or2_2 _17543_ (.A(_12630_),
    .B(_12626_),
    .X(_12631_));
 sky130_vsdinv _17544_ (.A(_12631_),
    .Y(_12632_));
 sky130_fd_sc_hd__a21oi_2 _17545_ (.A1(_12630_),
    .A2(_12626_),
    .B1(_12632_),
    .Y(_01583_));
 sky130_fd_sc_hd__o2bb2a_2 _17546_ (.A1_N(_02584_),
    .A2_N(\decoded_imm_uj[6] ),
    .B1(_12627_),
    .B2(_12628_),
    .X(_12633_));
 sky130_fd_sc_hd__nor2_2 _17547_ (.A(_02585_),
    .B(\decoded_imm_uj[7] ),
    .Y(_12634_));
 sky130_fd_sc_hd__a21o_2 _17548_ (.A1(_02585_),
    .A2(\decoded_imm_uj[7] ),
    .B1(_12634_),
    .X(_12635_));
 sky130_fd_sc_hd__o2bb2a_2 _17549_ (.A1_N(_12633_),
    .A2_N(_12635_),
    .B1(_12633_),
    .B2(_12635_),
    .X(_01584_));
 sky130_vsdinv _17550_ (.A(_02586_),
    .Y(_12636_));
 sky130_fd_sc_hd__or2_2 _17551_ (.A(_12636_),
    .B(_12631_),
    .X(_12637_));
 sky130_fd_sc_hd__o21a_2 _17552_ (.A1(_02586_),
    .A2(_12632_),
    .B1(_12637_),
    .X(_01587_));
 sky130_fd_sc_hd__o22a_2 _17553_ (.A1(_12630_),
    .A2(_12094_),
    .B1(_12633_),
    .B2(_12634_),
    .X(_12638_));
 sky130_fd_sc_hd__nor2_2 _17554_ (.A(_02586_),
    .B(\decoded_imm_uj[8] ),
    .Y(_12639_));
 sky130_fd_sc_hd__a21o_2 _17555_ (.A1(_02586_),
    .A2(\decoded_imm_uj[8] ),
    .B1(_12639_),
    .X(_12640_));
 sky130_fd_sc_hd__o2bb2a_2 _17556_ (.A1_N(_12638_),
    .A2_N(_12640_),
    .B1(_12638_),
    .B2(_12640_),
    .X(_01588_));
 sky130_vsdinv _17557_ (.A(_02587_),
    .Y(_12641_));
 sky130_fd_sc_hd__or2_2 _17558_ (.A(_12641_),
    .B(_12637_),
    .X(_12642_));
 sky130_vsdinv _17559_ (.A(_12642_),
    .Y(_12643_));
 sky130_fd_sc_hd__a21oi_2 _17560_ (.A1(_12641_),
    .A2(_12637_),
    .B1(_12643_),
    .Y(_01591_));
 sky130_fd_sc_hd__o22a_2 _17561_ (.A1(_12636_),
    .A2(_12098_),
    .B1(_12638_),
    .B2(_12639_),
    .X(_12644_));
 sky130_fd_sc_hd__nor2_2 _17562_ (.A(_02587_),
    .B(\decoded_imm_uj[9] ),
    .Y(_12645_));
 sky130_fd_sc_hd__a21o_2 _17563_ (.A1(_02587_),
    .A2(\decoded_imm_uj[9] ),
    .B1(_12645_),
    .X(_12646_));
 sky130_fd_sc_hd__o2bb2a_2 _17564_ (.A1_N(_12644_),
    .A2_N(_12646_),
    .B1(_12644_),
    .B2(_12646_),
    .X(_01592_));
 sky130_vsdinv _17565_ (.A(_02588_),
    .Y(_12647_));
 sky130_fd_sc_hd__or2_2 _17566_ (.A(_12647_),
    .B(_12642_),
    .X(_12648_));
 sky130_fd_sc_hd__o21a_2 _17567_ (.A1(_02588_),
    .A2(_12643_),
    .B1(_12648_),
    .X(_01595_));
 sky130_fd_sc_hd__o22a_2 _17568_ (.A1(_12641_),
    .A2(_12102_),
    .B1(_12644_),
    .B2(_12645_),
    .X(_12649_));
 sky130_fd_sc_hd__nor2_2 _17569_ (.A(_02588_),
    .B(\decoded_imm_uj[10] ),
    .Y(_12650_));
 sky130_fd_sc_hd__a21o_2 _17570_ (.A1(_02588_),
    .A2(\decoded_imm_uj[10] ),
    .B1(_12650_),
    .X(_12651_));
 sky130_fd_sc_hd__o2bb2a_2 _17571_ (.A1_N(_12649_),
    .A2_N(_12651_),
    .B1(_12649_),
    .B2(_12651_),
    .X(_01596_));
 sky130_vsdinv _17572_ (.A(_02589_),
    .Y(_12652_));
 sky130_fd_sc_hd__or2_2 _17573_ (.A(_12652_),
    .B(_12648_),
    .X(_12653_));
 sky130_vsdinv _17574_ (.A(_12653_),
    .Y(_12654_));
 sky130_fd_sc_hd__a21oi_2 _17575_ (.A1(_12652_),
    .A2(_12648_),
    .B1(_12654_),
    .Y(_01599_));
 sky130_fd_sc_hd__a22o_2 _17576_ (.A1(_02589_),
    .A2(\decoded_imm_uj[11] ),
    .B1(_12652_),
    .B2(_12112_),
    .X(_12655_));
 sky130_fd_sc_hd__o22a_2 _17577_ (.A1(_12647_),
    .A2(_12108_),
    .B1(_12649_),
    .B2(_12650_),
    .X(_12656_));
 sky130_fd_sc_hd__a2bb2oi_2 _17578_ (.A1_N(_12655_),
    .A2_N(_12656_),
    .B1(_12655_),
    .B2(_12656_),
    .Y(_01600_));
 sky130_vsdinv _17579_ (.A(_02561_),
    .Y(_12657_));
 sky130_fd_sc_hd__or2_2 _17580_ (.A(_12657_),
    .B(_12653_),
    .X(_12658_));
 sky130_fd_sc_hd__o21a_2 _17581_ (.A1(_02561_),
    .A2(_12654_),
    .B1(_12658_),
    .X(_01603_));
 sky130_fd_sc_hd__a22o_2 _17582_ (.A1(_02561_),
    .A2(\decoded_imm_uj[12] ),
    .B1(_12657_),
    .B2(_12116_),
    .X(_12659_));
 sky130_fd_sc_hd__o22a_2 _17583_ (.A1(_12652_),
    .A2(_12112_),
    .B1(_12655_),
    .B2(_12656_),
    .X(_12660_));
 sky130_fd_sc_hd__a2bb2oi_2 _17584_ (.A1_N(_12659_),
    .A2_N(_12660_),
    .B1(_12659_),
    .B2(_12660_),
    .Y(_01604_));
 sky130_vsdinv _17585_ (.A(_02562_),
    .Y(_12661_));
 sky130_fd_sc_hd__or2_2 _17586_ (.A(_12661_),
    .B(_12658_),
    .X(_12662_));
 sky130_vsdinv _17587_ (.A(_12662_),
    .Y(_12663_));
 sky130_fd_sc_hd__a21oi_2 _17588_ (.A1(_12661_),
    .A2(_12658_),
    .B1(_12663_),
    .Y(_01607_));
 sky130_fd_sc_hd__a22o_2 _17589_ (.A1(_02562_),
    .A2(\decoded_imm_uj[13] ),
    .B1(_12661_),
    .B2(_12123_),
    .X(_12664_));
 sky130_fd_sc_hd__o22a_2 _17590_ (.A1(_12657_),
    .A2(_12116_),
    .B1(_12659_),
    .B2(_12660_),
    .X(_12665_));
 sky130_fd_sc_hd__a2bb2oi_2 _17591_ (.A1_N(_12664_),
    .A2_N(_12665_),
    .B1(_12664_),
    .B2(_12665_),
    .Y(_01608_));
 sky130_vsdinv _17592_ (.A(_02563_),
    .Y(_12666_));
 sky130_fd_sc_hd__or2_2 _17593_ (.A(_12666_),
    .B(_12662_),
    .X(_12667_));
 sky130_fd_sc_hd__o21a_2 _17594_ (.A1(_02563_),
    .A2(_12663_),
    .B1(_12667_),
    .X(_01611_));
 sky130_fd_sc_hd__a22o_2 _17595_ (.A1(_02563_),
    .A2(\decoded_imm_uj[14] ),
    .B1(_12666_),
    .B2(_12127_),
    .X(_12668_));
 sky130_fd_sc_hd__o22a_2 _17596_ (.A1(_12661_),
    .A2(_12123_),
    .B1(_12664_),
    .B2(_12665_),
    .X(_12669_));
 sky130_fd_sc_hd__a2bb2oi_2 _17597_ (.A1_N(_12668_),
    .A2_N(_12669_),
    .B1(_12668_),
    .B2(_12669_),
    .Y(_01612_));
 sky130_vsdinv _17598_ (.A(_02564_),
    .Y(_12670_));
 sky130_fd_sc_hd__or2_2 _17599_ (.A(_12670_),
    .B(_12667_),
    .X(_12671_));
 sky130_vsdinv _17600_ (.A(_12671_),
    .Y(_12672_));
 sky130_fd_sc_hd__a21oi_2 _17601_ (.A1(_12670_),
    .A2(_12667_),
    .B1(_12672_),
    .Y(_01615_));
 sky130_fd_sc_hd__a22o_2 _17602_ (.A1(_02564_),
    .A2(\decoded_imm_uj[15] ),
    .B1(_12670_),
    .B2(_12130_),
    .X(_12673_));
 sky130_fd_sc_hd__o22a_2 _17603_ (.A1(_12666_),
    .A2(_12127_),
    .B1(_12668_),
    .B2(_12669_),
    .X(_12674_));
 sky130_fd_sc_hd__a2bb2oi_2 _17604_ (.A1_N(_12673_),
    .A2_N(_12674_),
    .B1(_12673_),
    .B2(_12674_),
    .Y(_01616_));
 sky130_vsdinv _17605_ (.A(_02565_),
    .Y(_12675_));
 sky130_fd_sc_hd__or2_2 _17606_ (.A(_12675_),
    .B(_12671_),
    .X(_12676_));
 sky130_fd_sc_hd__o21a_2 _17607_ (.A1(_02565_),
    .A2(_12672_),
    .B1(_12676_),
    .X(_01619_));
 sky130_fd_sc_hd__a22o_2 _17608_ (.A1(_02565_),
    .A2(\decoded_imm_uj[16] ),
    .B1(_12675_),
    .B2(_12135_),
    .X(_12677_));
 sky130_fd_sc_hd__o22a_2 _17609_ (.A1(_12670_),
    .A2(_12130_),
    .B1(_12673_),
    .B2(_12674_),
    .X(_12678_));
 sky130_fd_sc_hd__a2bb2oi_2 _17610_ (.A1_N(_12677_),
    .A2_N(_12678_),
    .B1(_12677_),
    .B2(_12678_),
    .Y(_01620_));
 sky130_vsdinv _17611_ (.A(_02566_),
    .Y(_12679_));
 sky130_fd_sc_hd__or2_2 _17612_ (.A(_12679_),
    .B(_12676_),
    .X(_12680_));
 sky130_vsdinv _17613_ (.A(_12680_),
    .Y(_12681_));
 sky130_fd_sc_hd__a21oi_2 _17614_ (.A1(_12679_),
    .A2(_12676_),
    .B1(_12681_),
    .Y(_01623_));
 sky130_fd_sc_hd__a22o_2 _17615_ (.A1(_02566_),
    .A2(\decoded_imm_uj[17] ),
    .B1(_12679_),
    .B2(_12139_),
    .X(_12682_));
 sky130_fd_sc_hd__o22a_2 _17616_ (.A1(_12675_),
    .A2(_12135_),
    .B1(_12677_),
    .B2(_12678_),
    .X(_12683_));
 sky130_fd_sc_hd__a2bb2oi_2 _17617_ (.A1_N(_12682_),
    .A2_N(_12683_),
    .B1(_12682_),
    .B2(_12683_),
    .Y(_01624_));
 sky130_vsdinv _17618_ (.A(_02567_),
    .Y(_12684_));
 sky130_fd_sc_hd__or2_2 _17619_ (.A(_12684_),
    .B(_12680_),
    .X(_12685_));
 sky130_fd_sc_hd__o21a_2 _17620_ (.A1(_02567_),
    .A2(_12681_),
    .B1(_12685_),
    .X(_01627_));
 sky130_fd_sc_hd__o22a_2 _17621_ (.A1(_12679_),
    .A2(_12139_),
    .B1(_12682_),
    .B2(_12683_),
    .X(_12686_));
 sky130_fd_sc_hd__nor2_2 _17622_ (.A(_02567_),
    .B(\decoded_imm_uj[18] ),
    .Y(_12687_));
 sky130_fd_sc_hd__a21o_2 _17623_ (.A1(_02567_),
    .A2(\decoded_imm_uj[18] ),
    .B1(_12687_),
    .X(_12688_));
 sky130_fd_sc_hd__o2bb2a_2 _17624_ (.A1_N(_12686_),
    .A2_N(_12688_),
    .B1(_12686_),
    .B2(_12688_),
    .X(_01628_));
 sky130_vsdinv _17625_ (.A(_02568_),
    .Y(_12689_));
 sky130_fd_sc_hd__or2_2 _17626_ (.A(_12689_),
    .B(_12685_),
    .X(_12690_));
 sky130_vsdinv _17627_ (.A(_12690_),
    .Y(_12691_));
 sky130_fd_sc_hd__a21oi_2 _17628_ (.A1(_12689_),
    .A2(_12685_),
    .B1(_12691_),
    .Y(_01631_));
 sky130_fd_sc_hd__a22o_2 _17629_ (.A1(_02568_),
    .A2(\decoded_imm_uj[19] ),
    .B1(_12689_),
    .B2(_12147_),
    .X(_12692_));
 sky130_fd_sc_hd__o22a_2 _17630_ (.A1(_12684_),
    .A2(_12143_),
    .B1(_12686_),
    .B2(_12687_),
    .X(_12693_));
 sky130_fd_sc_hd__a2bb2oi_2 _17631_ (.A1_N(_12692_),
    .A2_N(_12693_),
    .B1(_12692_),
    .B2(_12693_),
    .Y(_01632_));
 sky130_vsdinv _17632_ (.A(_02569_),
    .Y(_12694_));
 sky130_fd_sc_hd__or2_2 _17633_ (.A(_12694_),
    .B(_12690_),
    .X(_12695_));
 sky130_fd_sc_hd__o21a_2 _17634_ (.A1(_02569_),
    .A2(_12691_),
    .B1(_12695_),
    .X(_01635_));
 sky130_fd_sc_hd__o22a_2 _17635_ (.A1(_12689_),
    .A2(_12147_),
    .B1(_12692_),
    .B2(_12693_),
    .X(_12696_));
 sky130_fd_sc_hd__nor2_2 _17636_ (.A(_02569_),
    .B(\decoded_imm_uj[20] ),
    .Y(_12697_));
 sky130_fd_sc_hd__a21o_2 _17637_ (.A1(_02569_),
    .A2(_11707_),
    .B1(_12697_),
    .X(_12698_));
 sky130_fd_sc_hd__o2bb2a_2 _17638_ (.A1_N(_12696_),
    .A2_N(_12698_),
    .B1(_12696_),
    .B2(_12698_),
    .X(_01636_));
 sky130_vsdinv _17639_ (.A(_02570_),
    .Y(_12699_));
 sky130_fd_sc_hd__or2_2 _17640_ (.A(_12699_),
    .B(_12695_),
    .X(_12700_));
 sky130_vsdinv _17641_ (.A(_12700_),
    .Y(_12701_));
 sky130_fd_sc_hd__a21oi_2 _17642_ (.A1(_12699_),
    .A2(_12695_),
    .B1(_12701_),
    .Y(_01639_));
 sky130_fd_sc_hd__a22o_2 _17643_ (.A1(_02570_),
    .A2(_11705_),
    .B1(_12699_),
    .B2(_12155_),
    .X(_12702_));
 sky130_fd_sc_hd__o22a_2 _17644_ (.A1(_12694_),
    .A2(_12154_),
    .B1(_12696_),
    .B2(_12697_),
    .X(_12703_));
 sky130_fd_sc_hd__or2_2 _17645_ (.A(_12702_),
    .B(_12703_),
    .X(_12704_));
 sky130_fd_sc_hd__a21boi_2 _17646_ (.A1(_12702_),
    .A2(_12703_),
    .B1_N(_12704_),
    .Y(_01640_));
 sky130_vsdinv _17647_ (.A(_02572_),
    .Y(_12705_));
 sky130_fd_sc_hd__or2_2 _17648_ (.A(_12705_),
    .B(_12700_),
    .X(_12706_));
 sky130_fd_sc_hd__o21a_2 _17649_ (.A1(_02572_),
    .A2(_12701_),
    .B1(_12706_),
    .X(_01643_));
 sky130_fd_sc_hd__o22a_2 _17650_ (.A1(_12705_),
    .A2(_12155_),
    .B1(_02572_),
    .B2(_11705_),
    .X(_12707_));
 sky130_fd_sc_hd__o21ai_2 _17651_ (.A1(_12699_),
    .A2(_12158_),
    .B1(_12704_),
    .Y(_12708_));
 sky130_vsdinv _17652_ (.A(_12707_),
    .Y(_12709_));
 sky130_vsdinv _17653_ (.A(_12708_),
    .Y(_12710_));
 sky130_fd_sc_hd__o22a_2 _17654_ (.A1(_12707_),
    .A2(_12708_),
    .B1(_12709_),
    .B2(_12710_),
    .X(_01644_));
 sky130_vsdinv _17655_ (.A(_02573_),
    .Y(_12711_));
 sky130_fd_sc_hd__or2_2 _17656_ (.A(_12711_),
    .B(_12706_),
    .X(_12712_));
 sky130_vsdinv _17657_ (.A(_12712_),
    .Y(_12713_));
 sky130_fd_sc_hd__a21oi_2 _17658_ (.A1(_12711_),
    .A2(_12706_),
    .B1(_12713_),
    .Y(_01647_));
 sky130_fd_sc_hd__o22a_2 _17659_ (.A1(_12711_),
    .A2(_12155_),
    .B1(_02573_),
    .B2(_11705_),
    .X(_12714_));
 sky130_fd_sc_hd__or2_2 _17660_ (.A(_12704_),
    .B(_12709_),
    .X(_12715_));
 sky130_fd_sc_hd__o22a_2 _17661_ (.A1(_12699_),
    .A2(_12156_),
    .B1(_12705_),
    .B2(_12155_),
    .X(_12716_));
 sky130_fd_sc_hd__nand2_2 _17662_ (.A(_12715_),
    .B(_12716_),
    .Y(_12717_));
 sky130_fd_sc_hd__o2bb2a_2 _17663_ (.A1_N(_12714_),
    .A2_N(_12717_),
    .B1(_12714_),
    .B2(_12717_),
    .X(_01648_));
 sky130_vsdinv _17664_ (.A(_02574_),
    .Y(_12718_));
 sky130_fd_sc_hd__or2_2 _17665_ (.A(_12718_),
    .B(_12712_),
    .X(_12719_));
 sky130_fd_sc_hd__o21a_2 _17666_ (.A1(_02574_),
    .A2(_12713_),
    .B1(_12719_),
    .X(_01651_));
 sky130_fd_sc_hd__o22a_2 _17667_ (.A1(_12718_),
    .A2(_12155_),
    .B1(_02574_),
    .B2(_11705_),
    .X(_12720_));
 sky130_fd_sc_hd__a22o_2 _17668_ (.A1(_02573_),
    .A2(_11707_),
    .B1(_12714_),
    .B2(_12717_),
    .X(_12721_));
 sky130_vsdinv _17669_ (.A(_12720_),
    .Y(_12722_));
 sky130_vsdinv _17670_ (.A(_12721_),
    .Y(_12723_));
 sky130_fd_sc_hd__o22a_2 _17671_ (.A1(_12720_),
    .A2(_12721_),
    .B1(_12722_),
    .B2(_12723_),
    .X(_01652_));
 sky130_vsdinv _17672_ (.A(_02575_),
    .Y(_12724_));
 sky130_fd_sc_hd__or2_2 _17673_ (.A(_12724_),
    .B(_12719_),
    .X(_12725_));
 sky130_vsdinv _17674_ (.A(_12725_),
    .Y(_12726_));
 sky130_fd_sc_hd__a21oi_2 _17675_ (.A1(_12724_),
    .A2(_12719_),
    .B1(_12726_),
    .Y(_01655_));
 sky130_fd_sc_hd__a22o_2 _17676_ (.A1(_02575_),
    .A2(_11705_),
    .B1(_12724_),
    .B2(_12156_),
    .X(_12727_));
 sky130_vsdinv _17677_ (.A(_12714_),
    .Y(_12728_));
 sky130_fd_sc_hd__o22a_2 _17678_ (.A1(_12711_),
    .A2(_12156_),
    .B1(_12718_),
    .B2(_12156_),
    .X(_12729_));
 sky130_fd_sc_hd__o311a_2 _17679_ (.A1(_12728_),
    .A2(_12722_),
    .A3(_12715_),
    .B1(_12716_),
    .C1(_12729_),
    .X(_12730_));
 sky130_fd_sc_hd__or2_2 _17680_ (.A(_12727_),
    .B(_12730_),
    .X(_12731_));
 sky130_fd_sc_hd__a21boi_2 _17681_ (.A1(_12727_),
    .A2(_12730_),
    .B1_N(_12731_),
    .Y(_01656_));
 sky130_vsdinv _17682_ (.A(_02576_),
    .Y(_12732_));
 sky130_fd_sc_hd__or2_2 _17683_ (.A(_12732_),
    .B(_12725_),
    .X(_12733_));
 sky130_fd_sc_hd__o21a_2 _17684_ (.A1(_02576_),
    .A2(_12726_),
    .B1(_12733_),
    .X(_01659_));
 sky130_fd_sc_hd__o22a_2 _17685_ (.A1(_12732_),
    .A2(_12156_),
    .B1(_02576_),
    .B2(_11706_),
    .X(_12734_));
 sky130_fd_sc_hd__o21ai_2 _17686_ (.A1(_12724_),
    .A2(_12158_),
    .B1(_12731_),
    .Y(_12735_));
 sky130_vsdinv _17687_ (.A(_12734_),
    .Y(_12736_));
 sky130_vsdinv _17688_ (.A(_12735_),
    .Y(_12737_));
 sky130_fd_sc_hd__o22a_2 _17689_ (.A1(_12734_),
    .A2(_12735_),
    .B1(_12736_),
    .B2(_12737_),
    .X(_01660_));
 sky130_vsdinv _17690_ (.A(_02577_),
    .Y(_12738_));
 sky130_fd_sc_hd__or2_2 _17691_ (.A(_12738_),
    .B(_12733_),
    .X(_12739_));
 sky130_vsdinv _17692_ (.A(_12739_),
    .Y(_12740_));
 sky130_fd_sc_hd__a21oi_2 _17693_ (.A1(_12738_),
    .A2(_12733_),
    .B1(_12740_),
    .Y(_01663_));
 sky130_fd_sc_hd__o22a_2 _17694_ (.A1(_12738_),
    .A2(_12157_),
    .B1(_02577_),
    .B2(_11706_),
    .X(_12741_));
 sky130_fd_sc_hd__or2_2 _17695_ (.A(_12731_),
    .B(_12736_),
    .X(_12742_));
 sky130_fd_sc_hd__o22a_2 _17696_ (.A1(_12724_),
    .A2(_12157_),
    .B1(_12732_),
    .B2(_12157_),
    .X(_12743_));
 sky130_fd_sc_hd__nand2_2 _17697_ (.A(_12742_),
    .B(_12743_),
    .Y(_12744_));
 sky130_fd_sc_hd__o2bb2a_2 _17698_ (.A1_N(_12741_),
    .A2_N(_12744_),
    .B1(_12741_),
    .B2(_12744_),
    .X(_01664_));
 sky130_vsdinv _17699_ (.A(_02578_),
    .Y(_12745_));
 sky130_fd_sc_hd__or2_2 _17700_ (.A(_12745_),
    .B(_12739_),
    .X(_12746_));
 sky130_fd_sc_hd__o21a_2 _17701_ (.A1(_02578_),
    .A2(_12740_),
    .B1(_12746_),
    .X(_01667_));
 sky130_fd_sc_hd__o22a_2 _17702_ (.A1(_12745_),
    .A2(_12157_),
    .B1(_02578_),
    .B2(_11706_),
    .X(_12747_));
 sky130_fd_sc_hd__a22o_2 _17703_ (.A1(_02577_),
    .A2(_11706_),
    .B1(_12741_),
    .B2(_12744_),
    .X(_12748_));
 sky130_vsdinv _17704_ (.A(_12747_),
    .Y(_12749_));
 sky130_vsdinv _17705_ (.A(_12748_),
    .Y(_12750_));
 sky130_fd_sc_hd__o22a_2 _17706_ (.A1(_12747_),
    .A2(_12748_),
    .B1(_12749_),
    .B2(_12750_),
    .X(_01668_));
 sky130_vsdinv _17707_ (.A(_02579_),
    .Y(_12751_));
 sky130_fd_sc_hd__or2_2 _17708_ (.A(_12751_),
    .B(_12746_),
    .X(_12752_));
 sky130_vsdinv _17709_ (.A(_12752_),
    .Y(_12753_));
 sky130_fd_sc_hd__a21oi_2 _17710_ (.A1(_12751_),
    .A2(_12746_),
    .B1(_12753_),
    .Y(_01671_));
 sky130_fd_sc_hd__a22o_2 _17711_ (.A1(_02579_),
    .A2(_11706_),
    .B1(_12751_),
    .B2(_12158_),
    .X(_12754_));
 sky130_vsdinv _17712_ (.A(_12741_),
    .Y(_12755_));
 sky130_fd_sc_hd__o22a_2 _17713_ (.A1(_12738_),
    .A2(_12158_),
    .B1(_12745_),
    .B2(_12157_),
    .X(_12756_));
 sky130_fd_sc_hd__o311a_2 _17714_ (.A1(_12755_),
    .A2(_12749_),
    .A3(_12742_),
    .B1(_12743_),
    .C1(_12756_),
    .X(_12757_));
 sky130_fd_sc_hd__or2_2 _17715_ (.A(_12754_),
    .B(_12757_),
    .X(_12758_));
 sky130_vsdinv _17716_ (.A(_12758_),
    .Y(_12759_));
 sky130_fd_sc_hd__a21oi_2 _17717_ (.A1(_12754_),
    .A2(_12757_),
    .B1(_12759_),
    .Y(_01672_));
 sky130_vsdinv _17718_ (.A(_02580_),
    .Y(_12760_));
 sky130_fd_sc_hd__or2_2 _17719_ (.A(_12760_),
    .B(_12752_),
    .X(_12761_));
 sky130_fd_sc_hd__o21a_2 _17720_ (.A1(_02580_),
    .A2(_12753_),
    .B1(_12761_),
    .X(_01675_));
 sky130_fd_sc_hd__o22a_2 _17721_ (.A1(_02580_),
    .A2(_11707_),
    .B1(_12760_),
    .B2(_12174_),
    .X(_12762_));
 sky130_fd_sc_hd__o21ai_2 _17722_ (.A1(_12751_),
    .A2(_12174_),
    .B1(_12758_),
    .Y(_12763_));
 sky130_fd_sc_hd__a2bb2oi_2 _17723_ (.A1_N(_12762_),
    .A2_N(_12763_),
    .B1(_12762_),
    .B2(_12763_),
    .Y(_01676_));
 sky130_vsdinv _17724_ (.A(_02581_),
    .Y(_12764_));
 sky130_fd_sc_hd__a32o_2 _17725_ (.A1(_02580_),
    .A2(_12753_),
    .A3(_12764_),
    .B1(_02581_),
    .B2(_12761_),
    .X(_01679_));
 sky130_fd_sc_hd__o21ai_2 _17726_ (.A1(_02580_),
    .A2(_11707_),
    .B1(_12759_),
    .Y(_12765_));
 sky130_fd_sc_hd__o221ai_2 _17727_ (.A1(_12751_),
    .A2(_12174_),
    .B1(_12760_),
    .B2(_12174_),
    .C1(_12765_),
    .Y(_12766_));
 sky130_fd_sc_hd__a22o_2 _17728_ (.A1(_02581_),
    .A2(_12174_),
    .B1(_12764_),
    .B2(_11707_),
    .X(_12767_));
 sky130_fd_sc_hd__a2bb2oi_2 _17729_ (.A1_N(_12766_),
    .A2_N(_12767_),
    .B1(_12766_),
    .B2(_12767_),
    .Y(_01680_));
 sky130_fd_sc_hd__or2_2 _17730_ (.A(\mem_wordsize[2] ),
    .B(\mem_wordsize[1] ),
    .X(_12768_));
 sky130_vsdinv _17731_ (.A(_12768_),
    .Y(_12769_));
 sky130_fd_sc_hd__buf_1 _17732_ (.A(_12769_),
    .X(_01683_));
 sky130_fd_sc_hd__buf_1 _17733_ (.A(_12451_),
    .X(_12770_));
 sky130_fd_sc_hd__a211o_2 _17734_ (.A1(_12770_),
    .A2(\mem_wordsize[2] ),
    .B1(_12769_),
    .C1(_00304_),
    .X(mem_la_wstrb[0]));
 sky130_fd_sc_hd__and2_2 _17735_ (.A(mem_la_write),
    .B(mem_la_wstrb[0]),
    .X(_01684_));
 sky130_fd_sc_hd__and3_2 _17736_ (.A(_10811_),
    .B(_00301_),
    .C(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__buf_1 _17737_ (.A(_12768_),
    .X(_12771_));
 sky130_fd_sc_hd__or2_2 _17738_ (.A(_11862_),
    .B(_12196_),
    .X(_12772_));
 sky130_fd_sc_hd__o211a_2 _17739_ (.A1(_11862_),
    .A2(_12359_),
    .B1(_12771_),
    .C1(_12772_),
    .X(_12773_));
 sky130_fd_sc_hd__nor2_2 _17740_ (.A(_11396_),
    .B(_12773_),
    .Y(_01687_));
 sky130_fd_sc_hd__and3_2 _17741_ (.A(_10811_),
    .B(_00301_),
    .C(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__or2_2 _17742_ (.A(_12770_),
    .B(_11863_),
    .X(_12774_));
 sky130_fd_sc_hd__buf_1 _17743_ (.A(_12774_),
    .X(_12775_));
 sky130_fd_sc_hd__o211a_2 _17744_ (.A1(_12770_),
    .A2(_12359_),
    .B1(_12771_),
    .C1(_12775_),
    .X(_12776_));
 sky130_fd_sc_hd__nor2_2 _17745_ (.A(_11396_),
    .B(_12776_),
    .Y(_01690_));
 sky130_fd_sc_hd__and3_2 _17746_ (.A(_10811_),
    .B(_00301_),
    .C(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__or2_2 _17747_ (.A(_12770_),
    .B(_12196_),
    .X(_12777_));
 sky130_fd_sc_hd__o211a_2 _17748_ (.A1(_12770_),
    .A2(_12207_),
    .B1(_12768_),
    .C1(_12777_),
    .X(_12778_));
 sky130_fd_sc_hd__nor2_2 _17749_ (.A(_11396_),
    .B(_12778_),
    .Y(_01693_));
 sky130_fd_sc_hd__and3_2 _17750_ (.A(_10811_),
    .B(_00301_),
    .C(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__or2_2 _17751_ (.A(\irq_pending[1] ),
    .B(irq[1]),
    .X(_12779_));
 sky130_fd_sc_hd__buf_1 _17752_ (.A(_12779_),
    .X(_01697_));
 sky130_fd_sc_hd__inv_2 _17753_ (.A(_01697_),
    .Y(_01696_));
 sky130_fd_sc_hd__nor2_2 _17754_ (.A(_10510_),
    .B(_01696_),
    .Y(_01698_));
 sky130_fd_sc_hd__and3_2 _17755_ (.A(_11251_),
    .B(_00297_),
    .C(_12178_),
    .X(_12780_));
 sky130_fd_sc_hd__nand2_2 _17756_ (.A(_12182_),
    .B(_12780_),
    .Y(_02217_));
 sky130_vsdinv _17757_ (.A(_02217_),
    .Y(_01700_));
 sky130_fd_sc_hd__o21a_2 _17758_ (.A1(irq_active),
    .A2(\irq_mask[1] ),
    .B1(_01696_),
    .X(_01701_));
 sky130_fd_sc_hd__o22ai_2 _17759_ (.A1(_01696_),
    .A2(_12780_),
    .B1(_12182_),
    .B2(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__buf_1 _17760_ (.A(_10459_),
    .X(_12781_));
 sky130_fd_sc_hd__and2_2 _17761_ (.A(_12781_),
    .B(_00354_),
    .X(_01706_));
 sky130_vsdinv _17762_ (.A(mem_rdata[0]),
    .Y(_01707_));
 sky130_vsdinv _17763_ (.A(mem_rdata[24]),
    .Y(_12782_));
 sky130_fd_sc_hd__buf_1 _17764_ (.A(_12777_),
    .X(_12783_));
 sky130_vsdinv _17765_ (.A(mem_rdata[8]),
    .Y(_01812_));
 sky130_fd_sc_hd__buf_1 _17766_ (.A(_12772_),
    .X(_12784_));
 sky130_vsdinv _17767_ (.A(mem_rdata[16]),
    .Y(_12785_));
 sky130_fd_sc_hd__or2_2 _17768_ (.A(_12785_),
    .B(_12775_),
    .X(_12786_));
 sky130_fd_sc_hd__o221a_2 _17769_ (.A1(_12782_),
    .A2(_12783_),
    .B1(_01812_),
    .B2(_12784_),
    .C1(_12786_),
    .X(_01708_));
 sky130_vsdinv _17770_ (.A(_01710_),
    .Y(_12787_));
 sky130_fd_sc_hd__o22a_2 _17771_ (.A1(_12373_),
    .A2(_01709_),
    .B1(_12360_),
    .B2(_12787_),
    .X(_01711_));
 sky130_fd_sc_hd__buf_1 _17772_ (.A(_11766_),
    .X(_12788_));
 sky130_fd_sc_hd__buf_1 _17773_ (.A(_11773_),
    .X(_12789_));
 sky130_fd_sc_hd__or2_2 _17774_ (.A(_10909_),
    .B(_11768_),
    .X(_12790_));
 sky130_fd_sc_hd__o221a_2 _17775_ (.A1(_10877_),
    .A2(_12788_),
    .B1(_12789_),
    .B2(_11148_),
    .C1(_12790_),
    .X(_01715_));
 sky130_fd_sc_hd__buf_1 _17776_ (.A(_11735_),
    .X(_12791_));
 sky130_fd_sc_hd__buf_1 _17777_ (.A(_11741_),
    .X(_12792_));
 sky130_fd_sc_hd__o21ai_2 _17778_ (.A1(instr_setq),
    .A2(instr_getq),
    .B1(\cpuregs_rs1[0] ),
    .Y(_12793_));
 sky130_fd_sc_hd__o221a_2 _17779_ (.A1(_12791_),
    .A2(_12409_),
    .B1(_11079_),
    .B2(_12792_),
    .C1(_12793_),
    .X(_01718_));
 sky130_fd_sc_hd__buf_1 _17780_ (.A(_11030_),
    .X(_12794_));
 sky130_fd_sc_hd__o2bb2a_2 _17781_ (.A1_N(_11085_),
    .A2_N(_01713_),
    .B1(_12794_),
    .B2(_01719_),
    .X(_12795_));
 sky130_fd_sc_hd__buf_1 _17782_ (.A(_10609_),
    .X(_12796_));
 sky130_fd_sc_hd__a221o_2 _17783_ (.A1(\decoded_imm[0] ),
    .A2(\reg_next_pc[0] ),
    .B1(_11715_),
    .B2(_12447_),
    .C1(_12796_),
    .X(_12797_));
 sky130_fd_sc_hd__o211ai_2 _17784_ (.A1(_12256_),
    .A2(_01712_),
    .B1(_12795_),
    .C1(_12797_),
    .Y(_01720_));
 sky130_vsdinv _17785_ (.A(mem_rdata[1]),
    .Y(_01721_));
 sky130_vsdinv _17786_ (.A(mem_rdata[25]),
    .Y(_12798_));
 sky130_vsdinv _17787_ (.A(mem_rdata[9]),
    .Y(_01826_));
 sky130_vsdinv _17788_ (.A(mem_rdata[17]),
    .Y(_12799_));
 sky130_fd_sc_hd__or2_2 _17789_ (.A(_12799_),
    .B(_12775_),
    .X(_12800_));
 sky130_fd_sc_hd__o221a_2 _17790_ (.A1(_12798_),
    .A2(_12783_),
    .B1(_01826_),
    .B2(_12784_),
    .C1(_12800_),
    .X(_01722_));
 sky130_vsdinv _17791_ (.A(_01724_),
    .Y(_12801_));
 sky130_fd_sc_hd__o22a_2 _17792_ (.A1(_12373_),
    .A2(_01723_),
    .B1(_12360_),
    .B2(_12801_),
    .X(_01725_));
 sky130_fd_sc_hd__or2_2 _17793_ (.A(_10876_),
    .B(_11766_),
    .X(_12802_));
 sky130_fd_sc_hd__o221a_2 _17794_ (.A1(_10908_),
    .A2(_11768_),
    .B1(_12789_),
    .B2(_11147_),
    .C1(_12802_),
    .X(_01729_));
 sky130_fd_sc_hd__buf_1 _17795_ (.A(_10620_),
    .X(_12803_));
 sky130_fd_sc_hd__buf_1 _17796_ (.A(_12803_),
    .X(_12804_));
 sky130_fd_sc_hd__nand2_2 _17797_ (.A(_12804_),
    .B(\cpuregs_rs1[1] ),
    .Y(_12805_));
 sky130_fd_sc_hd__o221a_2 _17798_ (.A1(_12791_),
    .A2(_12408_),
    .B1(_10510_),
    .B2(_12792_),
    .C1(_12805_),
    .X(_01731_));
 sky130_fd_sc_hd__a22o_2 _17799_ (.A1(\reg_pc[1] ),
    .A2(\decoded_imm[1] ),
    .B1(_12449_),
    .B2(_12058_),
    .X(_12806_));
 sky130_fd_sc_hd__or3_2 _17800_ (.A(_11715_),
    .B(_12447_),
    .C(_12806_),
    .X(_12807_));
 sky130_fd_sc_hd__o21ai_2 _17801_ (.A1(_11715_),
    .A2(_12447_),
    .B1(_12806_),
    .Y(_12808_));
 sky130_fd_sc_hd__buf_1 _17802_ (.A(_10459_),
    .X(_12809_));
 sky130_fd_sc_hd__buf_1 _17803_ (.A(_10639_),
    .X(_12810_));
 sky130_fd_sc_hd__o2bb2a_2 _17804_ (.A1_N(_12810_),
    .A2_N(_01727_),
    .B1(_11080_),
    .B2(_01732_),
    .X(_12811_));
 sky130_fd_sc_hd__o21ai_2 _17805_ (.A1(_12809_),
    .A2(_01726_),
    .B1(_12811_),
    .Y(_12812_));
 sky130_fd_sc_hd__a31o_2 _17806_ (.A1(_12364_),
    .A2(_12807_),
    .A3(_12808_),
    .B1(_12812_),
    .X(_01733_));
 sky130_vsdinv _17807_ (.A(mem_rdata[2]),
    .Y(_01734_));
 sky130_vsdinv _17808_ (.A(mem_rdata[26]),
    .Y(_12813_));
 sky130_vsdinv _17809_ (.A(mem_rdata[10]),
    .Y(_01839_));
 sky130_vsdinv _17810_ (.A(mem_rdata[18]),
    .Y(_12814_));
 sky130_fd_sc_hd__or2_2 _17811_ (.A(_12814_),
    .B(_12775_),
    .X(_12815_));
 sky130_fd_sc_hd__o221a_2 _17812_ (.A1(_12813_),
    .A2(_12783_),
    .B1(_01839_),
    .B2(_12784_),
    .C1(_12815_),
    .X(_01735_));
 sky130_vsdinv _17813_ (.A(_01737_),
    .Y(_12816_));
 sky130_fd_sc_hd__o22a_2 _17814_ (.A1(_12373_),
    .A2(_01736_),
    .B1(_12360_),
    .B2(_12816_),
    .X(_01738_));
 sky130_fd_sc_hd__or2_2 _17815_ (.A(_10907_),
    .B(_11768_),
    .X(_12817_));
 sky130_fd_sc_hd__o221a_2 _17816_ (.A1(_10875_),
    .A2(_12788_),
    .B1(_12789_),
    .B2(_11146_),
    .C1(_12817_),
    .X(_01742_));
 sky130_vsdinv _17817_ (.A(\timer[2] ),
    .Y(_12818_));
 sky130_fd_sc_hd__nand2_2 _17818_ (.A(_12804_),
    .B(\cpuregs_rs1[2] ),
    .Y(_12819_));
 sky130_fd_sc_hd__o221a_2 _17819_ (.A1(_12791_),
    .A2(_12818_),
    .B1(_10511_),
    .B2(_12792_),
    .C1(_12819_),
    .X(_01744_));
 sky130_fd_sc_hd__o2bb2a_2 _17820_ (.A1_N(_11085_),
    .A2_N(_01740_),
    .B1(_12794_),
    .B2(_01745_),
    .X(_12820_));
 sky130_fd_sc_hd__o21ai_2 _17821_ (.A1(_12449_),
    .A2(_12058_),
    .B1(_12807_),
    .Y(_12821_));
 sky130_fd_sc_hd__nor2_2 _17822_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .Y(_12822_));
 sky130_fd_sc_hd__a21oi_2 _17823_ (.A1(\reg_pc[2] ),
    .A2(\decoded_imm[2] ),
    .B1(_12822_),
    .Y(_12823_));
 sky130_vsdinv _17824_ (.A(_12821_),
    .Y(_12824_));
 sky130_vsdinv _17825_ (.A(_12823_),
    .Y(_12825_));
 sky130_fd_sc_hd__a221o_2 _17826_ (.A1(_12821_),
    .A2(_12823_),
    .B1(_12824_),
    .B2(_12825_),
    .C1(_10610_),
    .X(_12826_));
 sky130_fd_sc_hd__o211ai_2 _17827_ (.A1(_12256_),
    .A2(_01739_),
    .B1(_12820_),
    .C1(_12826_),
    .Y(_01746_));
 sky130_vsdinv _17828_ (.A(mem_rdata[3]),
    .Y(_01747_));
 sky130_vsdinv _17829_ (.A(mem_rdata[27]),
    .Y(_12827_));
 sky130_vsdinv _17830_ (.A(mem_rdata[11]),
    .Y(_01852_));
 sky130_vsdinv _17831_ (.A(mem_rdata[19]),
    .Y(_12828_));
 sky130_fd_sc_hd__or2_2 _17832_ (.A(_12828_),
    .B(_12775_),
    .X(_12829_));
 sky130_fd_sc_hd__o221a_2 _17833_ (.A1(_12827_),
    .A2(_12783_),
    .B1(_01852_),
    .B2(_12784_),
    .C1(_12829_),
    .X(_01748_));
 sky130_vsdinv _17834_ (.A(_01750_),
    .Y(_12830_));
 sky130_fd_sc_hd__o22a_2 _17835_ (.A1(_12373_),
    .A2(_01749_),
    .B1(_12360_),
    .B2(_12830_),
    .X(_01751_));
 sky130_fd_sc_hd__or2_2 _17836_ (.A(_10906_),
    .B(_11768_),
    .X(_12831_));
 sky130_fd_sc_hd__o221a_2 _17837_ (.A1(_10874_),
    .A2(_12788_),
    .B1(_12789_),
    .B2(_11145_),
    .C1(_12831_),
    .X(_01755_));
 sky130_fd_sc_hd__buf_1 _17838_ (.A(_12803_),
    .X(_12832_));
 sky130_fd_sc_hd__buf_1 _17839_ (.A(instr_timer),
    .X(_12833_));
 sky130_fd_sc_hd__buf_1 _17840_ (.A(_12833_),
    .X(_12834_));
 sky130_fd_sc_hd__buf_1 _17841_ (.A(instr_maskirq),
    .X(_12835_));
 sky130_fd_sc_hd__buf_1 _17842_ (.A(_12835_),
    .X(_12836_));
 sky130_fd_sc_hd__a22o_2 _17843_ (.A1(_12834_),
    .A2(\timer[3] ),
    .B1(\irq_mask[3] ),
    .B2(_12836_),
    .X(_12837_));
 sky130_fd_sc_hd__a21oi_2 _17844_ (.A1(_12832_),
    .A2(\cpuregs_rs1[3] ),
    .B1(_12837_),
    .Y(_01757_));
 sky130_fd_sc_hd__o2bb2a_2 _17845_ (.A1_N(_11085_),
    .A2_N(_01753_),
    .B1(_11031_),
    .B2(_01758_),
    .X(_12838_));
 sky130_fd_sc_hd__o22a_2 _17846_ (.A1(_02073_),
    .A2(_12065_),
    .B1(_12824_),
    .B2(_12822_),
    .X(_12839_));
 sky130_vsdinv _17847_ (.A(_12839_),
    .Y(_12840_));
 sky130_fd_sc_hd__nor2_2 _17848_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .Y(_12841_));
 sky130_fd_sc_hd__a21oi_2 _17849_ (.A1(\reg_pc[3] ),
    .A2(\decoded_imm[3] ),
    .B1(_12841_),
    .Y(_12842_));
 sky130_vsdinv _17850_ (.A(_12842_),
    .Y(_12843_));
 sky130_fd_sc_hd__a221o_2 _17851_ (.A1(_12840_),
    .A2(_12842_),
    .B1(_12839_),
    .B2(_12843_),
    .C1(_10610_),
    .X(_12844_));
 sky130_fd_sc_hd__o211ai_2 _17852_ (.A1(_12256_),
    .A2(_01752_),
    .B1(_12838_),
    .C1(_12844_),
    .Y(_01759_));
 sky130_vsdinv _17853_ (.A(mem_rdata[4]),
    .Y(_01760_));
 sky130_vsdinv _17854_ (.A(mem_rdata[28]),
    .Y(_12845_));
 sky130_vsdinv _17855_ (.A(mem_rdata[12]),
    .Y(_01865_));
 sky130_vsdinv _17856_ (.A(mem_rdata[20]),
    .Y(_12846_));
 sky130_fd_sc_hd__or2_2 _17857_ (.A(_12846_),
    .B(_12775_),
    .X(_12847_));
 sky130_fd_sc_hd__o221a_2 _17858_ (.A1(_12845_),
    .A2(_12783_),
    .B1(_01865_),
    .B2(_12784_),
    .C1(_12847_),
    .X(_01761_));
 sky130_vsdinv _17859_ (.A(_01763_),
    .Y(_12848_));
 sky130_fd_sc_hd__o22a_2 _17860_ (.A1(_12373_),
    .A2(_01762_),
    .B1(_12360_),
    .B2(_12848_),
    .X(_01764_));
 sky130_fd_sc_hd__or2_2 _17861_ (.A(_10905_),
    .B(_11768_),
    .X(_12849_));
 sky130_fd_sc_hd__o221a_2 _17862_ (.A1(_10873_),
    .A2(_12788_),
    .B1(_12789_),
    .B2(_11144_),
    .C1(_12849_),
    .X(_01768_));
 sky130_fd_sc_hd__a22o_2 _17863_ (.A1(_12834_),
    .A2(\timer[4] ),
    .B1(\irq_mask[4] ),
    .B2(_12836_),
    .X(_12850_));
 sky130_fd_sc_hd__a21oi_2 _17864_ (.A1(_12832_),
    .A2(\cpuregs_rs1[4] ),
    .B1(_12850_),
    .Y(_01770_));
 sky130_fd_sc_hd__o22ai_2 _17865_ (.A1(_12458_),
    .A2(_12071_),
    .B1(_12839_),
    .B2(_12841_),
    .Y(_12851_));
 sky130_fd_sc_hd__o22a_2 _17866_ (.A1(_12463_),
    .A2(_12077_),
    .B1(\reg_pc[4] ),
    .B2(\decoded_imm[4] ),
    .X(_12852_));
 sky130_fd_sc_hd__or2_2 _17867_ (.A(_12851_),
    .B(_12852_),
    .X(_12853_));
 sky130_fd_sc_hd__nand2_2 _17868_ (.A(_12851_),
    .B(_12852_),
    .Y(_12854_));
 sky130_fd_sc_hd__o2bb2a_2 _17869_ (.A1_N(_12810_),
    .A2_N(_01766_),
    .B1(_11080_),
    .B2(_01771_),
    .X(_12855_));
 sky130_fd_sc_hd__o21ai_2 _17870_ (.A1(_12809_),
    .A2(_01765_),
    .B1(_12855_),
    .Y(_12856_));
 sky130_fd_sc_hd__a31o_2 _17871_ (.A1(_12364_),
    .A2(_12853_),
    .A3(_12854_),
    .B1(_12856_),
    .X(_01772_));
 sky130_vsdinv _17872_ (.A(mem_rdata[5]),
    .Y(_01773_));
 sky130_vsdinv _17873_ (.A(mem_rdata[29]),
    .Y(_12857_));
 sky130_vsdinv _17874_ (.A(mem_rdata[13]),
    .Y(_01878_));
 sky130_vsdinv _17875_ (.A(mem_rdata[21]),
    .Y(_12858_));
 sky130_fd_sc_hd__or2_2 _17876_ (.A(_12858_),
    .B(_12774_),
    .X(_12859_));
 sky130_fd_sc_hd__o221a_2 _17877_ (.A1(_12857_),
    .A2(_12783_),
    .B1(_01878_),
    .B2(_12784_),
    .C1(_12859_),
    .X(_01774_));
 sky130_vsdinv _17878_ (.A(_01776_),
    .Y(_12860_));
 sky130_fd_sc_hd__o22a_2 _17879_ (.A1(_12372_),
    .A2(_01775_),
    .B1(_12359_),
    .B2(_12860_),
    .X(_01777_));
 sky130_fd_sc_hd__buf_1 _17880_ (.A(_10617_),
    .X(_12861_));
 sky130_fd_sc_hd__buf_1 _17881_ (.A(_12861_),
    .X(_12862_));
 sky130_fd_sc_hd__or2_2 _17882_ (.A(_10904_),
    .B(_12862_),
    .X(_12863_));
 sky130_fd_sc_hd__o221a_2 _17883_ (.A1(_10872_),
    .A2(_12788_),
    .B1(_12789_),
    .B2(_11143_),
    .C1(_12863_),
    .X(_01781_));
 sky130_fd_sc_hd__buf_1 _17884_ (.A(_12803_),
    .X(_12864_));
 sky130_fd_sc_hd__nand2_2 _17885_ (.A(_12864_),
    .B(\cpuregs_rs1[5] ),
    .Y(_12865_));
 sky130_fd_sc_hd__o221a_2 _17886_ (.A1(_12791_),
    .A2(_12411_),
    .B1(_10528_),
    .B2(_12792_),
    .C1(_12865_),
    .X(_01783_));
 sky130_fd_sc_hd__buf_1 _17887_ (.A(_12810_),
    .X(_12866_));
 sky130_fd_sc_hd__nor2_2 _17888_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .Y(_12867_));
 sky130_fd_sc_hd__a21oi_2 _17889_ (.A1(\reg_pc[5] ),
    .A2(\decoded_imm[5] ),
    .B1(_12867_),
    .Y(_12868_));
 sky130_fd_sc_hd__o21ai_2 _17890_ (.A1(_12463_),
    .A2(_12077_),
    .B1(_12854_),
    .Y(_12869_));
 sky130_fd_sc_hd__or2_2 _17891_ (.A(_12868_),
    .B(_12869_),
    .X(_12870_));
 sky130_fd_sc_hd__a21oi_2 _17892_ (.A1(_12868_),
    .A2(_12869_),
    .B1(_12274_),
    .Y(_12871_));
 sky130_fd_sc_hd__o22ai_2 _17893_ (.A1(_12255_),
    .A2(_01778_),
    .B1(_12369_),
    .B2(_01784_),
    .Y(_12872_));
 sky130_fd_sc_hd__a221o_2 _17894_ (.A1(_12866_),
    .A2(_01779_),
    .B1(_12870_),
    .B2(_12871_),
    .C1(_12872_),
    .X(_01785_));
 sky130_vsdinv _17895_ (.A(mem_rdata[6]),
    .Y(_01786_));
 sky130_vsdinv _17896_ (.A(mem_rdata[30]),
    .Y(_12873_));
 sky130_vsdinv _17897_ (.A(mem_rdata[14]),
    .Y(_01891_));
 sky130_vsdinv _17898_ (.A(mem_rdata[22]),
    .Y(_12874_));
 sky130_fd_sc_hd__or2_2 _17899_ (.A(_12874_),
    .B(_12774_),
    .X(_12875_));
 sky130_fd_sc_hd__o221a_2 _17900_ (.A1(_12873_),
    .A2(_12777_),
    .B1(_01891_),
    .B2(_12772_),
    .C1(_12875_),
    .X(_01787_));
 sky130_vsdinv _17901_ (.A(_01789_),
    .Y(_12876_));
 sky130_fd_sc_hd__o22a_2 _17902_ (.A1(_12372_),
    .A2(_01788_),
    .B1(_12359_),
    .B2(_12876_),
    .X(_01790_));
 sky130_fd_sc_hd__buf_1 _17903_ (.A(_11773_),
    .X(_12877_));
 sky130_fd_sc_hd__or2_2 _17904_ (.A(_10903_),
    .B(_12862_),
    .X(_12878_));
 sky130_fd_sc_hd__o221a_2 _17905_ (.A1(_10871_),
    .A2(_12788_),
    .B1(_12877_),
    .B2(_11142_),
    .C1(_12878_),
    .X(_01794_));
 sky130_fd_sc_hd__a22o_2 _17906_ (.A1(_12834_),
    .A2(\timer[6] ),
    .B1(\irq_mask[6] ),
    .B2(_12836_),
    .X(_12879_));
 sky130_fd_sc_hd__a21oi_2 _17907_ (.A1(_12832_),
    .A2(\cpuregs_rs1[6] ),
    .B1(_12879_),
    .Y(_01796_));
 sky130_fd_sc_hd__o32a_2 _17908_ (.A1(_12463_),
    .A2(_12077_),
    .A3(_12867_),
    .B1(_12468_),
    .B2(_12084_),
    .X(_12880_));
 sky130_vsdinv _17909_ (.A(_12880_),
    .Y(_12881_));
 sky130_fd_sc_hd__a31o_2 _17910_ (.A1(_12852_),
    .A2(_12868_),
    .A3(_12851_),
    .B1(_12881_),
    .X(_12882_));
 sky130_fd_sc_hd__o22a_2 _17911_ (.A1(_12473_),
    .A2(_12091_),
    .B1(\reg_pc[6] ),
    .B2(\decoded_imm[6] ),
    .X(_12883_));
 sky130_fd_sc_hd__or2_2 _17912_ (.A(_12882_),
    .B(_12883_),
    .X(_12884_));
 sky130_fd_sc_hd__nand2_2 _17913_ (.A(_12882_),
    .B(_12883_),
    .Y(_12885_));
 sky130_fd_sc_hd__o2bb2a_2 _17914_ (.A1_N(_12810_),
    .A2_N(_01792_),
    .B1(_11080_),
    .B2(_01797_),
    .X(_12886_));
 sky130_fd_sc_hd__o21ai_2 _17915_ (.A1(_12809_),
    .A2(_01791_),
    .B1(_12886_),
    .Y(_12887_));
 sky130_fd_sc_hd__a31o_2 _17916_ (.A1(_12364_),
    .A2(_12884_),
    .A3(_12885_),
    .B1(_12887_),
    .X(_01798_));
 sky130_vsdinv _17917_ (.A(mem_rdata[7]),
    .Y(_01799_));
 sky130_vsdinv _17918_ (.A(mem_rdata[31]),
    .Y(_12888_));
 sky130_vsdinv _17919_ (.A(mem_rdata[15]),
    .Y(_01904_));
 sky130_vsdinv _17920_ (.A(mem_rdata[23]),
    .Y(_12889_));
 sky130_fd_sc_hd__or2_2 _17921_ (.A(_12889_),
    .B(_12774_),
    .X(_12890_));
 sky130_fd_sc_hd__o221a_2 _17922_ (.A1(_12888_),
    .A2(_12777_),
    .B1(_01904_),
    .B2(_12772_),
    .C1(_12890_),
    .X(_01800_));
 sky130_vsdinv _17923_ (.A(_01802_),
    .Y(_12891_));
 sky130_fd_sc_hd__o22a_2 _17924_ (.A1(_12372_),
    .A2(_01801_),
    .B1(_12359_),
    .B2(_12891_),
    .X(_01803_));
 sky130_fd_sc_hd__buf_1 _17925_ (.A(_11766_),
    .X(_12892_));
 sky130_fd_sc_hd__or2_2 _17926_ (.A(_10902_),
    .B(_12862_),
    .X(_12893_));
 sky130_fd_sc_hd__o221a_2 _17927_ (.A1(_10870_),
    .A2(_12892_),
    .B1(_12877_),
    .B2(_11141_),
    .C1(_12893_),
    .X(_01807_));
 sky130_fd_sc_hd__nand2_2 _17928_ (.A(_12864_),
    .B(\cpuregs_rs1[7] ),
    .Y(_12894_));
 sky130_fd_sc_hd__o221a_2 _17929_ (.A1(_12791_),
    .A2(_12413_),
    .B1(_10529_),
    .B2(_12792_),
    .C1(_12894_),
    .X(_01809_));
 sky130_fd_sc_hd__nor2_2 _17930_ (.A(\reg_pc[7] ),
    .B(\decoded_imm[7] ),
    .Y(_12895_));
 sky130_fd_sc_hd__a21oi_2 _17931_ (.A1(\reg_pc[7] ),
    .A2(\decoded_imm[7] ),
    .B1(_12895_),
    .Y(_12896_));
 sky130_fd_sc_hd__o21ai_2 _17932_ (.A1(_12473_),
    .A2(_12091_),
    .B1(_12885_),
    .Y(_12897_));
 sky130_fd_sc_hd__or2_2 _17933_ (.A(_12896_),
    .B(_12897_),
    .X(_12898_));
 sky130_fd_sc_hd__a21oi_2 _17934_ (.A1(_12896_),
    .A2(_12897_),
    .B1(_12796_),
    .Y(_12899_));
 sky130_fd_sc_hd__o22ai_2 _17935_ (.A1(_12794_),
    .A2(_01810_),
    .B1(_12781_),
    .B2(_01804_),
    .Y(_12900_));
 sky130_fd_sc_hd__a221o_2 _17936_ (.A1(_12866_),
    .A2(_01805_),
    .B1(_12898_),
    .B2(_12899_),
    .C1(_12900_),
    .X(_01811_));
 sky130_fd_sc_hd__buf_1 _17937_ (.A(\mem_wordsize[2] ),
    .X(_12901_));
 sky130_fd_sc_hd__buf_1 _17938_ (.A(_12901_),
    .X(_12902_));
 sky130_fd_sc_hd__nand2_2 _17939_ (.A(_12902_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_2 _17940_ (.A(latched_is_lb),
    .B(latched_is_lh),
    .Y(_01816_));
 sky130_vsdinv _17941_ (.A(latched_is_lb),
    .Y(_12903_));
 sky130_fd_sc_hd__buf_1 _17942_ (.A(_12903_),
    .X(_12904_));
 sky130_fd_sc_hd__buf_1 _17943_ (.A(_01804_),
    .X(_12905_));
 sky130_vsdinv _17944_ (.A(latched_is_lh),
    .Y(_12906_));
 sky130_fd_sc_hd__buf_1 _17945_ (.A(_12906_),
    .X(_12907_));
 sky130_fd_sc_hd__o22a_2 _17946_ (.A1(_12904_),
    .A2(_12905_),
    .B1(_12907_),
    .B2(_01815_),
    .X(_01817_));
 sky130_fd_sc_hd__or2_2 _17947_ (.A(_10901_),
    .B(_12862_),
    .X(_12908_));
 sky130_fd_sc_hd__o221a_2 _17948_ (.A1(_10869_),
    .A2(_12892_),
    .B1(_12877_),
    .B2(_11140_),
    .C1(_12908_),
    .X(_01821_));
 sky130_fd_sc_hd__a22o_2 _17949_ (.A1(_12834_),
    .A2(\timer[8] ),
    .B1(\irq_mask[8] ),
    .B2(_12836_),
    .X(_12909_));
 sky130_fd_sc_hd__a21oi_2 _17950_ (.A1(_12832_),
    .A2(\cpuregs_rs1[8] ),
    .B1(_12909_),
    .Y(_01823_));
 sky130_fd_sc_hd__o32a_2 _17951_ (.A1(_12473_),
    .A2(_12090_),
    .A3(_12895_),
    .B1(_12478_),
    .B2(_12093_),
    .X(_12910_));
 sky130_vsdinv _17952_ (.A(_12910_),
    .Y(_12911_));
 sky130_fd_sc_hd__a31o_2 _17953_ (.A1(_12883_),
    .A2(_12896_),
    .A3(_12882_),
    .B1(_12911_),
    .X(_12912_));
 sky130_fd_sc_hd__o22a_2 _17954_ (.A1(_12483_),
    .A2(_12096_),
    .B1(\reg_pc[8] ),
    .B2(\decoded_imm[8] ),
    .X(_12913_));
 sky130_fd_sc_hd__or2_2 _17955_ (.A(_12912_),
    .B(_12913_),
    .X(_12914_));
 sky130_fd_sc_hd__nand2_2 _17956_ (.A(_12912_),
    .B(_12913_),
    .Y(_12915_));
 sky130_fd_sc_hd__o2bb2a_2 _17957_ (.A1_N(_12810_),
    .A2_N(_01819_),
    .B1(_11080_),
    .B2(_01824_),
    .X(_12916_));
 sky130_fd_sc_hd__o21ai_2 _17958_ (.A1(_12809_),
    .A2(_01818_),
    .B1(_12916_),
    .Y(_12917_));
 sky130_fd_sc_hd__a31o_2 _17959_ (.A1(_12364_),
    .A2(_12914_),
    .A3(_12915_),
    .B1(_12917_),
    .X(_01825_));
 sky130_fd_sc_hd__nand2_2 _17960_ (.A(_12902_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__o22a_2 _17961_ (.A1(_12904_),
    .A2(_12905_),
    .B1(_12907_),
    .B2(_01829_),
    .X(_01830_));
 sky130_fd_sc_hd__or2_2 _17962_ (.A(_10900_),
    .B(_12862_),
    .X(_12918_));
 sky130_fd_sc_hd__o221a_2 _17963_ (.A1(_10868_),
    .A2(_12892_),
    .B1(_12877_),
    .B2(_11139_),
    .C1(_12918_),
    .X(_01834_));
 sky130_fd_sc_hd__nand2_2 _17964_ (.A(_12864_),
    .B(\cpuregs_rs1[9] ),
    .Y(_12919_));
 sky130_fd_sc_hd__o221a_2 _17965_ (.A1(_12791_),
    .A2(_12415_),
    .B1(_10547_),
    .B2(_12792_),
    .C1(_12919_),
    .X(_01836_));
 sky130_fd_sc_hd__nor2_2 _17966_ (.A(\reg_pc[9] ),
    .B(\decoded_imm[9] ),
    .Y(_12920_));
 sky130_fd_sc_hd__a21oi_2 _17967_ (.A1(\reg_pc[9] ),
    .A2(\decoded_imm[9] ),
    .B1(_12920_),
    .Y(_12921_));
 sky130_fd_sc_hd__o21ai_2 _17968_ (.A1(_12483_),
    .A2(_12097_),
    .B1(_12915_),
    .Y(_12922_));
 sky130_fd_sc_hd__or2_2 _17969_ (.A(_12921_),
    .B(_12922_),
    .X(_12923_));
 sky130_fd_sc_hd__a21oi_2 _17970_ (.A1(_12921_),
    .A2(_12922_),
    .B1(_12796_),
    .Y(_12924_));
 sky130_fd_sc_hd__o22ai_2 _17971_ (.A1(_12255_),
    .A2(_01831_),
    .B1(_12369_),
    .B2(_01837_),
    .Y(_12925_));
 sky130_fd_sc_hd__a221o_2 _17972_ (.A1(_12866_),
    .A2(_01832_),
    .B1(_12923_),
    .B2(_12924_),
    .C1(_12925_),
    .X(_01838_));
 sky130_fd_sc_hd__nand2_2 _17973_ (.A(_12902_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__o22a_2 _17974_ (.A1(_12904_),
    .A2(_12905_),
    .B1(_12907_),
    .B2(_01842_),
    .X(_01843_));
 sky130_fd_sc_hd__or2_2 _17975_ (.A(_10899_),
    .B(_12862_),
    .X(_12926_));
 sky130_fd_sc_hd__o221a_2 _17976_ (.A1(_10867_),
    .A2(_12892_),
    .B1(_12877_),
    .B2(_11138_),
    .C1(_12926_),
    .X(_01847_));
 sky130_fd_sc_hd__a22o_2 _17977_ (.A1(_12834_),
    .A2(\timer[10] ),
    .B1(\irq_mask[10] ),
    .B2(_12836_),
    .X(_12927_));
 sky130_fd_sc_hd__a21oi_2 _17978_ (.A1(_12832_),
    .A2(\cpuregs_rs1[10] ),
    .B1(_12927_),
    .Y(_01849_));
 sky130_fd_sc_hd__o22a_2 _17979_ (.A1(_12496_),
    .A2(_12105_),
    .B1(\reg_pc[10] ),
    .B2(\decoded_imm[10] ),
    .X(_12928_));
 sky130_fd_sc_hd__o32a_2 _17980_ (.A1(_12483_),
    .A2(_12096_),
    .A3(_12920_),
    .B1(_12492_),
    .B2(_12101_),
    .X(_12929_));
 sky130_vsdinv _17981_ (.A(_12929_),
    .Y(_12930_));
 sky130_fd_sc_hd__a31o_2 _17982_ (.A1(_12913_),
    .A2(_12921_),
    .A3(_12912_),
    .B1(_12930_),
    .X(_12931_));
 sky130_fd_sc_hd__or2_2 _17983_ (.A(_12928_),
    .B(_12931_),
    .X(_12932_));
 sky130_fd_sc_hd__nand2_2 _17984_ (.A(_12928_),
    .B(_12931_),
    .Y(_12933_));
 sky130_fd_sc_hd__buf_1 _17985_ (.A(_10469_),
    .X(_12934_));
 sky130_fd_sc_hd__o2bb2a_2 _17986_ (.A1_N(_12810_),
    .A2_N(_01845_),
    .B1(_12934_),
    .B2(_01850_),
    .X(_12935_));
 sky130_fd_sc_hd__o21ai_2 _17987_ (.A1(_12809_),
    .A2(_01844_),
    .B1(_12935_),
    .Y(_12936_));
 sky130_fd_sc_hd__a31o_2 _17988_ (.A1(_12364_),
    .A2(_12932_),
    .A3(_12933_),
    .B1(_12936_),
    .X(_01851_));
 sky130_fd_sc_hd__nand2_2 _17989_ (.A(_12902_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__o22a_2 _17990_ (.A1(_12904_),
    .A2(_12905_),
    .B1(_12907_),
    .B2(_01855_),
    .X(_01856_));
 sky130_fd_sc_hd__buf_1 _17991_ (.A(_12861_),
    .X(_12937_));
 sky130_fd_sc_hd__or2_2 _17992_ (.A(_10898_),
    .B(_12937_),
    .X(_12938_));
 sky130_fd_sc_hd__o221a_2 _17993_ (.A1(_10866_),
    .A2(_12892_),
    .B1(_12877_),
    .B2(_11137_),
    .C1(_12938_),
    .X(_01860_));
 sky130_fd_sc_hd__buf_1 _17994_ (.A(_11734_),
    .X(_12939_));
 sky130_fd_sc_hd__buf_1 _17995_ (.A(_10678_),
    .X(_12940_));
 sky130_fd_sc_hd__nand2_2 _17996_ (.A(_12864_),
    .B(\cpuregs_rs1[11] ),
    .Y(_12941_));
 sky130_fd_sc_hd__o221a_2 _17997_ (.A1(_12939_),
    .A2(_12417_),
    .B1(_10548_),
    .B2(_12940_),
    .C1(_12941_),
    .X(_01862_));
 sky130_fd_sc_hd__buf_1 _17998_ (.A(_10603_),
    .X(_04073_));
 sky130_fd_sc_hd__o22a_2 _17999_ (.A1(_12502_),
    .A2(_12111_),
    .B1(\reg_pc[11] ),
    .B2(\decoded_imm[11] ),
    .X(_04074_));
 sky130_fd_sc_hd__o21ai_2 _18000_ (.A1(_12496_),
    .A2(_12105_),
    .B1(_12933_),
    .Y(_04075_));
 sky130_fd_sc_hd__nand2_2 _18001_ (.A(_04074_),
    .B(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__or2_2 _18002_ (.A(_04074_),
    .B(_04075_),
    .X(_04077_));
 sky130_fd_sc_hd__buf_1 _18003_ (.A(_10459_),
    .X(_04078_));
 sky130_fd_sc_hd__buf_1 _18004_ (.A(_11084_),
    .X(_04079_));
 sky130_fd_sc_hd__o2bb2a_2 _18005_ (.A1_N(_04079_),
    .A2_N(_01858_),
    .B1(_12934_),
    .B2(_01863_),
    .X(_04080_));
 sky130_fd_sc_hd__o21ai_2 _18006_ (.A1(_04078_),
    .A2(_01857_),
    .B1(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__a31o_2 _18007_ (.A1(_04073_),
    .A2(_04076_),
    .A3(_04077_),
    .B1(_04081_),
    .X(_01864_));
 sky130_fd_sc_hd__nand2_2 _18008_ (.A(_12902_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__o22a_2 _18009_ (.A1(_12904_),
    .A2(_12905_),
    .B1(_12907_),
    .B2(_01868_),
    .X(_01869_));
 sky130_fd_sc_hd__buf_1 _18010_ (.A(_11773_),
    .X(_04082_));
 sky130_fd_sc_hd__or2_2 _18011_ (.A(_10897_),
    .B(_12937_),
    .X(_04083_));
 sky130_fd_sc_hd__o221a_2 _18012_ (.A1(_10865_),
    .A2(_12892_),
    .B1(_04082_),
    .B2(_11136_),
    .C1(_04083_),
    .X(_01873_));
 sky130_fd_sc_hd__a22o_2 _18013_ (.A1(_12834_),
    .A2(\timer[12] ),
    .B1(\irq_mask[12] ),
    .B2(_12836_),
    .X(_04084_));
 sky130_fd_sc_hd__a21oi_2 _18014_ (.A1(_12832_),
    .A2(\cpuregs_rs1[12] ),
    .B1(_04084_),
    .Y(_01875_));
 sky130_fd_sc_hd__o22a_2 _18015_ (.A1(_12506_),
    .A2(_12115_),
    .B1(\reg_pc[12] ),
    .B2(\decoded_imm[12] ),
    .X(_04085_));
 sky130_fd_sc_hd__o21ai_2 _18016_ (.A1(_12502_),
    .A2(_12111_),
    .B1(_04076_),
    .Y(_04086_));
 sky130_fd_sc_hd__or2_2 _18017_ (.A(_04085_),
    .B(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__nand2_2 _18018_ (.A(_04085_),
    .B(_04086_),
    .Y(_04088_));
 sky130_fd_sc_hd__o2bb2a_2 _18019_ (.A1_N(_04079_),
    .A2_N(_01871_),
    .B1(_12934_),
    .B2(_01876_),
    .X(_04089_));
 sky130_fd_sc_hd__o21ai_2 _18020_ (.A1(_04078_),
    .A2(_01870_),
    .B1(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__a31o_2 _18021_ (.A1(_04073_),
    .A2(_04087_),
    .A3(_04088_),
    .B1(_04090_),
    .X(_01877_));
 sky130_fd_sc_hd__nand2_2 _18022_ (.A(_12902_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__o22a_2 _18023_ (.A1(_12904_),
    .A2(_12905_),
    .B1(_12907_),
    .B2(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__buf_1 _18024_ (.A(_11766_),
    .X(_04091_));
 sky130_fd_sc_hd__or2_2 _18025_ (.A(_10896_),
    .B(_12937_),
    .X(_04092_));
 sky130_fd_sc_hd__o221a_2 _18026_ (.A1(_10864_),
    .A2(_04091_),
    .B1(_04082_),
    .B2(_11135_),
    .C1(_04092_),
    .X(_01886_));
 sky130_fd_sc_hd__nand2_2 _18027_ (.A(_12864_),
    .B(\cpuregs_rs1[13] ),
    .Y(_04093_));
 sky130_fd_sc_hd__o221a_2 _18028_ (.A1(_12939_),
    .A2(_12419_),
    .B1(_10535_),
    .B2(_12940_),
    .C1(_04093_),
    .X(_01888_));
 sky130_fd_sc_hd__o22a_2 _18029_ (.A1(_12510_),
    .A2(_12122_),
    .B1(\reg_pc[13] ),
    .B2(\decoded_imm[13] ),
    .X(_04094_));
 sky130_fd_sc_hd__o21ai_2 _18030_ (.A1(_12506_),
    .A2(_12115_),
    .B1(_04088_),
    .Y(_04095_));
 sky130_fd_sc_hd__nand2_2 _18031_ (.A(_04094_),
    .B(_04095_),
    .Y(_04096_));
 sky130_fd_sc_hd__or2_2 _18032_ (.A(_04094_),
    .B(_04095_),
    .X(_04097_));
 sky130_fd_sc_hd__o2bb2a_2 _18033_ (.A1_N(_04079_),
    .A2_N(_01884_),
    .B1(_12934_),
    .B2(_01889_),
    .X(_04098_));
 sky130_fd_sc_hd__o21ai_2 _18034_ (.A1(_04078_),
    .A2(_01883_),
    .B1(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__a31o_2 _18035_ (.A1(_04073_),
    .A2(_04096_),
    .A3(_04097_),
    .B1(_04099_),
    .X(_01890_));
 sky130_fd_sc_hd__buf_1 _18036_ (.A(_12901_),
    .X(_04100_));
 sky130_fd_sc_hd__nand2_2 _18037_ (.A(_04100_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__o22a_2 _18038_ (.A1(_12903_),
    .A2(_01804_),
    .B1(_12906_),
    .B2(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__or2_2 _18039_ (.A(_10895_),
    .B(_12937_),
    .X(_04101_));
 sky130_fd_sc_hd__o221a_2 _18040_ (.A1(_10863_),
    .A2(_04091_),
    .B1(_04082_),
    .B2(_11134_),
    .C1(_04101_),
    .X(_01899_));
 sky130_fd_sc_hd__buf_1 _18041_ (.A(_12803_),
    .X(_04102_));
 sky130_fd_sc_hd__buf_1 _18042_ (.A(_12833_),
    .X(_04103_));
 sky130_fd_sc_hd__buf_1 _18043_ (.A(_12835_),
    .X(_04104_));
 sky130_fd_sc_hd__a22o_2 _18044_ (.A1(_04103_),
    .A2(\timer[14] ),
    .B1(\irq_mask[14] ),
    .B2(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__a21oi_2 _18045_ (.A1(_04102_),
    .A2(\cpuregs_rs1[14] ),
    .B1(_04105_),
    .Y(_01901_));
 sky130_fd_sc_hd__o22a_2 _18046_ (.A1(_12515_),
    .A2(_12126_),
    .B1(\reg_pc[14] ),
    .B2(\decoded_imm[14] ),
    .X(_04106_));
 sky130_fd_sc_hd__o21ai_2 _18047_ (.A1(_12510_),
    .A2(_12122_),
    .B1(_04096_),
    .Y(_04107_));
 sky130_fd_sc_hd__or2_2 _18048_ (.A(_04106_),
    .B(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__nand2_2 _18049_ (.A(_04106_),
    .B(_04107_),
    .Y(_04109_));
 sky130_fd_sc_hd__o2bb2a_2 _18050_ (.A1_N(_04079_),
    .A2_N(_01897_),
    .B1(_12934_),
    .B2(_01902_),
    .X(_04110_));
 sky130_fd_sc_hd__o21ai_2 _18051_ (.A1(_04078_),
    .A2(_01896_),
    .B1(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__a31o_2 _18052_ (.A1(_04073_),
    .A2(_04108_),
    .A3(_04109_),
    .B1(_04111_),
    .X(_01903_));
 sky130_fd_sc_hd__nand2_2 _18053_ (.A(_04100_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__o22a_2 _18054_ (.A1(_12903_),
    .A2(_01804_),
    .B1(_12906_),
    .B2(_01907_),
    .X(_01908_));
 sky130_fd_sc_hd__or2_2 _18055_ (.A(_10894_),
    .B(_12937_),
    .X(_04112_));
 sky130_fd_sc_hd__o221a_2 _18056_ (.A1(_10862_),
    .A2(_04091_),
    .B1(_04082_),
    .B2(_11133_),
    .C1(_04112_),
    .X(_01912_));
 sky130_fd_sc_hd__nand2_2 _18057_ (.A(_12864_),
    .B(\cpuregs_rs1[15] ),
    .Y(_04113_));
 sky130_fd_sc_hd__o221a_2 _18058_ (.A1(_12939_),
    .A2(_12421_),
    .B1(_10536_),
    .B2(_12940_),
    .C1(_04113_),
    .X(_01914_));
 sky130_fd_sc_hd__o22a_2 _18059_ (.A1(_12519_),
    .A2(_12129_),
    .B1(\reg_pc[15] ),
    .B2(\decoded_imm[15] ),
    .X(_04114_));
 sky130_fd_sc_hd__o21ai_2 _18060_ (.A1(_12515_),
    .A2(_12126_),
    .B1(_04109_),
    .Y(_04115_));
 sky130_fd_sc_hd__nand2_2 _18061_ (.A(_04114_),
    .B(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__or2_2 _18062_ (.A(_04114_),
    .B(_04115_),
    .X(_04117_));
 sky130_fd_sc_hd__o2bb2a_2 _18063_ (.A1_N(_04079_),
    .A2_N(_01910_),
    .B1(_12934_),
    .B2(_01915_),
    .X(_04118_));
 sky130_fd_sc_hd__o21ai_2 _18064_ (.A1(_04078_),
    .A2(_01909_),
    .B1(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__a31o_2 _18065_ (.A1(_04073_),
    .A2(_04116_),
    .A3(_04117_),
    .B1(_04119_),
    .X(_01916_));
 sky130_fd_sc_hd__buf_1 _18066_ (.A(_12768_),
    .X(_04120_));
 sky130_fd_sc_hd__or2_2 _18067_ (.A(_12785_),
    .B(_04120_),
    .X(_01917_));
 sky130_fd_sc_hd__or2_2 _18068_ (.A(_10893_),
    .B(_12937_),
    .X(_04121_));
 sky130_fd_sc_hd__o221a_2 _18069_ (.A1(_10861_),
    .A2(_04091_),
    .B1(_04082_),
    .B2(_11132_),
    .C1(_04121_),
    .X(_01921_));
 sky130_fd_sc_hd__a22o_2 _18070_ (.A1(_04103_),
    .A2(\timer[16] ),
    .B1(\irq_mask[16] ),
    .B2(_04104_),
    .X(_04122_));
 sky130_fd_sc_hd__a21oi_2 _18071_ (.A1(_04102_),
    .A2(\cpuregs_rs1[16] ),
    .B1(_04122_),
    .Y(_01923_));
 sky130_fd_sc_hd__o21ai_2 _18072_ (.A1(_12519_),
    .A2(_12129_),
    .B1(_04116_),
    .Y(_04123_));
 sky130_fd_sc_hd__o22a_2 _18073_ (.A1(_12523_),
    .A2(_12133_),
    .B1(\reg_pc[16] ),
    .B2(\decoded_imm[16] ),
    .X(_04124_));
 sky130_fd_sc_hd__or2_2 _18074_ (.A(_04123_),
    .B(_04124_),
    .X(_04125_));
 sky130_fd_sc_hd__nand2_2 _18075_ (.A(_04123_),
    .B(_04124_),
    .Y(_04126_));
 sky130_fd_sc_hd__buf_1 _18076_ (.A(_10469_),
    .X(_04127_));
 sky130_fd_sc_hd__o2bb2a_2 _18077_ (.A1_N(_04079_),
    .A2_N(_01919_),
    .B1(_04127_),
    .B2(_01924_),
    .X(_04128_));
 sky130_fd_sc_hd__o21ai_2 _18078_ (.A1(_04078_),
    .A2(_01918_),
    .B1(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__a31o_2 _18079_ (.A1(_04073_),
    .A2(_04125_),
    .A3(_04126_),
    .B1(_04129_),
    .X(_01925_));
 sky130_fd_sc_hd__or2_2 _18080_ (.A(_12799_),
    .B(_04120_),
    .X(_01926_));
 sky130_fd_sc_hd__buf_1 _18081_ (.A(_12861_),
    .X(_04130_));
 sky130_fd_sc_hd__or2_2 _18082_ (.A(_10892_),
    .B(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__o221a_2 _18083_ (.A1(_10860_),
    .A2(_04091_),
    .B1(_04082_),
    .B2(_11131_),
    .C1(_04131_),
    .X(_01930_));
 sky130_fd_sc_hd__a22o_2 _18084_ (.A1(_04103_),
    .A2(\timer[17] ),
    .B1(\irq_mask[17] ),
    .B2(_04104_),
    .X(_04132_));
 sky130_fd_sc_hd__a21oi_2 _18085_ (.A1(_04102_),
    .A2(\cpuregs_rs1[17] ),
    .B1(_04132_),
    .Y(_01932_));
 sky130_fd_sc_hd__nor2_2 _18086_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .Y(_04133_));
 sky130_fd_sc_hd__a21oi_2 _18087_ (.A1(\reg_pc[17] ),
    .A2(\decoded_imm[17] ),
    .B1(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__o21ai_2 _18088_ (.A1(_12523_),
    .A2(_12134_),
    .B1(_04126_),
    .Y(_04135_));
 sky130_fd_sc_hd__or2_2 _18089_ (.A(_04134_),
    .B(_04135_),
    .X(_04136_));
 sky130_fd_sc_hd__a21oi_2 _18090_ (.A1(_04134_),
    .A2(_04135_),
    .B1(_12796_),
    .Y(_04137_));
 sky130_fd_sc_hd__o22ai_2 _18091_ (.A1(_12255_),
    .A2(_01927_),
    .B1(_12794_),
    .B2(_01933_),
    .Y(_04138_));
 sky130_fd_sc_hd__a221o_2 _18092_ (.A1(_12866_),
    .A2(_01928_),
    .B1(_04136_),
    .B2(_04137_),
    .C1(_04138_),
    .X(_01934_));
 sky130_fd_sc_hd__or2_2 _18093_ (.A(_12814_),
    .B(_04120_),
    .X(_01935_));
 sky130_fd_sc_hd__buf_1 _18094_ (.A(_10618_),
    .X(_04139_));
 sky130_fd_sc_hd__or2_2 _18095_ (.A(_10891_),
    .B(_04130_),
    .X(_04140_));
 sky130_fd_sc_hd__o221a_2 _18096_ (.A1(_10859_),
    .A2(_04091_),
    .B1(_04139_),
    .B2(_11130_),
    .C1(_04140_),
    .X(_01939_));
 sky130_fd_sc_hd__buf_1 _18097_ (.A(_12803_),
    .X(_04141_));
 sky130_fd_sc_hd__nand2_2 _18098_ (.A(_04141_),
    .B(\cpuregs_rs1[18] ),
    .Y(_04142_));
 sky130_fd_sc_hd__o221a_2 _18099_ (.A1(_12939_),
    .A2(_12378_),
    .B1(_11052_),
    .B2(_12940_),
    .C1(_04142_),
    .X(_01941_));
 sky130_fd_sc_hd__buf_1 _18100_ (.A(_10603_),
    .X(_04143_));
 sky130_fd_sc_hd__o22a_2 _18101_ (.A1(_12533_),
    .A2(_12142_),
    .B1(\reg_pc[18] ),
    .B2(\decoded_imm[18] ),
    .X(_04144_));
 sky130_fd_sc_hd__o32a_2 _18102_ (.A1(_12523_),
    .A2(_12133_),
    .A3(_04133_),
    .B1(_12529_),
    .B2(_12138_),
    .X(_04145_));
 sky130_vsdinv _18103_ (.A(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__a31o_2 _18104_ (.A1(_04124_),
    .A2(_04134_),
    .A3(_04123_),
    .B1(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__or2_2 _18105_ (.A(_04144_),
    .B(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__nand2_2 _18106_ (.A(_04144_),
    .B(_04147_),
    .Y(_04149_));
 sky130_fd_sc_hd__buf_1 _18107_ (.A(_10459_),
    .X(_04150_));
 sky130_fd_sc_hd__buf_1 _18108_ (.A(_10639_),
    .X(_04151_));
 sky130_fd_sc_hd__o2bb2a_2 _18109_ (.A1_N(_04151_),
    .A2_N(_01937_),
    .B1(_04127_),
    .B2(_01942_),
    .X(_04152_));
 sky130_fd_sc_hd__o21ai_2 _18110_ (.A1(_04150_),
    .A2(_01936_),
    .B1(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__a31o_2 _18111_ (.A1(_04143_),
    .A2(_04148_),
    .A3(_04149_),
    .B1(_04153_),
    .X(_01943_));
 sky130_fd_sc_hd__or2_2 _18112_ (.A(_12828_),
    .B(_04120_),
    .X(_01944_));
 sky130_fd_sc_hd__buf_1 _18113_ (.A(_10616_),
    .X(_04154_));
 sky130_fd_sc_hd__or2_2 _18114_ (.A(_10890_),
    .B(_04130_),
    .X(_04155_));
 sky130_fd_sc_hd__o221a_2 _18115_ (.A1(_10858_),
    .A2(_04154_),
    .B1(_04139_),
    .B2(_11129_),
    .C1(_04155_),
    .X(_01948_));
 sky130_fd_sc_hd__a22o_2 _18116_ (.A1(_04103_),
    .A2(\timer[19] ),
    .B1(\irq_mask[19] ),
    .B2(_04104_),
    .X(_04156_));
 sky130_fd_sc_hd__a21oi_2 _18117_ (.A1(_04102_),
    .A2(\cpuregs_rs1[19] ),
    .B1(_04156_),
    .Y(_01950_));
 sky130_fd_sc_hd__o22a_2 _18118_ (.A1(_12539_),
    .A2(_12146_),
    .B1(\reg_pc[19] ),
    .B2(\decoded_imm[19] ),
    .X(_04157_));
 sky130_fd_sc_hd__o21ai_2 _18119_ (.A1(_12533_),
    .A2(_12142_),
    .B1(_04149_),
    .Y(_04158_));
 sky130_fd_sc_hd__nand2_2 _18120_ (.A(_04157_),
    .B(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__or2_2 _18121_ (.A(_04157_),
    .B(_04158_),
    .X(_04160_));
 sky130_fd_sc_hd__o2bb2a_2 _18122_ (.A1_N(_04151_),
    .A2_N(_01946_),
    .B1(_04127_),
    .B2(_01951_),
    .X(_04161_));
 sky130_fd_sc_hd__o21ai_2 _18123_ (.A1(_04150_),
    .A2(_01945_),
    .B1(_04161_),
    .Y(_04162_));
 sky130_fd_sc_hd__a31o_2 _18124_ (.A1(_04143_),
    .A2(_04159_),
    .A3(_04160_),
    .B1(_04162_),
    .X(_01952_));
 sky130_fd_sc_hd__or2_2 _18125_ (.A(_12846_),
    .B(_04120_),
    .X(_01953_));
 sky130_fd_sc_hd__or2_2 _18126_ (.A(_10889_),
    .B(_04130_),
    .X(_04163_));
 sky130_fd_sc_hd__o221a_2 _18127_ (.A1(_10857_),
    .A2(_04154_),
    .B1(_04139_),
    .B2(_11128_),
    .C1(_04163_),
    .X(_01957_));
 sky130_fd_sc_hd__nand2_2 _18128_ (.A(_04141_),
    .B(\cpuregs_rs1[20] ),
    .Y(_04164_));
 sky130_fd_sc_hd__o221a_2 _18129_ (.A1(_12939_),
    .A2(_12423_),
    .B1(_10553_),
    .B2(_12940_),
    .C1(_04164_),
    .X(_01959_));
 sky130_fd_sc_hd__o22a_2 _18130_ (.A1(_12544_),
    .A2(_12435_),
    .B1(\reg_pc[20] ),
    .B2(\decoded_imm[20] ),
    .X(_04165_));
 sky130_fd_sc_hd__o21ai_2 _18131_ (.A1(_12539_),
    .A2(_12146_),
    .B1(_04159_),
    .Y(_04166_));
 sky130_fd_sc_hd__or2_2 _18132_ (.A(_04165_),
    .B(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__nand2_2 _18133_ (.A(_04165_),
    .B(_04166_),
    .Y(_04168_));
 sky130_fd_sc_hd__o2bb2a_2 _18134_ (.A1_N(_04151_),
    .A2_N(_01955_),
    .B1(_04127_),
    .B2(_01960_),
    .X(_04169_));
 sky130_fd_sc_hd__o21ai_2 _18135_ (.A1(_04150_),
    .A2(_01954_),
    .B1(_04169_),
    .Y(_04170_));
 sky130_fd_sc_hd__a31o_2 _18136_ (.A1(_04143_),
    .A2(_04167_),
    .A3(_04168_),
    .B1(_04170_),
    .X(_01961_));
 sky130_fd_sc_hd__or2_2 _18137_ (.A(_12858_),
    .B(_04120_),
    .X(_01962_));
 sky130_fd_sc_hd__or2_2 _18138_ (.A(_10888_),
    .B(_04130_),
    .X(_04171_));
 sky130_fd_sc_hd__o221a_2 _18139_ (.A1(_10856_),
    .A2(_04154_),
    .B1(_04139_),
    .B2(_11127_),
    .C1(_04171_),
    .X(_01966_));
 sky130_fd_sc_hd__a22o_2 _18140_ (.A1(_04103_),
    .A2(\timer[21] ),
    .B1(\irq_mask[21] ),
    .B2(_04104_),
    .X(_04172_));
 sky130_fd_sc_hd__a21oi_2 _18141_ (.A1(_04102_),
    .A2(\cpuregs_rs1[21] ),
    .B1(_04172_),
    .Y(_01968_));
 sky130_fd_sc_hd__o22a_2 _18142_ (.A1(_12548_),
    .A2(_12436_),
    .B1(\reg_pc[21] ),
    .B2(\decoded_imm[21] ),
    .X(_04173_));
 sky130_fd_sc_hd__o21ai_2 _18143_ (.A1(_12544_),
    .A2(_12435_),
    .B1(_04168_),
    .Y(_04174_));
 sky130_fd_sc_hd__nand2_2 _18144_ (.A(_04173_),
    .B(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__or2_2 _18145_ (.A(_04173_),
    .B(_04174_),
    .X(_04176_));
 sky130_fd_sc_hd__o2bb2a_2 _18146_ (.A1_N(_04151_),
    .A2_N(_01964_),
    .B1(_04127_),
    .B2(_01969_),
    .X(_04177_));
 sky130_fd_sc_hd__o21ai_2 _18147_ (.A1(_04150_),
    .A2(_01963_),
    .B1(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__a31o_2 _18148_ (.A1(_04143_),
    .A2(_04175_),
    .A3(_04176_),
    .B1(_04178_),
    .X(_01970_));
 sky130_fd_sc_hd__buf_1 _18149_ (.A(_12768_),
    .X(_04179_));
 sky130_fd_sc_hd__or2_2 _18150_ (.A(_12874_),
    .B(_04179_),
    .X(_01971_));
 sky130_fd_sc_hd__or2_2 _18151_ (.A(_10887_),
    .B(_04130_),
    .X(_04180_));
 sky130_fd_sc_hd__o221a_2 _18152_ (.A1(_10855_),
    .A2(_04154_),
    .B1(_04139_),
    .B2(_11126_),
    .C1(_04180_),
    .X(_01975_));
 sky130_fd_sc_hd__nand2_2 _18153_ (.A(_04141_),
    .B(\cpuregs_rs1[22] ),
    .Y(_04181_));
 sky130_fd_sc_hd__o221a_2 _18154_ (.A1(_12939_),
    .A2(_12425_),
    .B1(_10554_),
    .B2(_12940_),
    .C1(_04181_),
    .X(_01977_));
 sky130_fd_sc_hd__o22a_2 _18155_ (.A1(_12552_),
    .A2(_12438_),
    .B1(\reg_pc[22] ),
    .B2(\decoded_imm[22] ),
    .X(_04182_));
 sky130_fd_sc_hd__o21ai_2 _18156_ (.A1(_12548_),
    .A2(_12436_),
    .B1(_04175_),
    .Y(_04183_));
 sky130_fd_sc_hd__or2_2 _18157_ (.A(_04182_),
    .B(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__nand2_2 _18158_ (.A(_04182_),
    .B(_04183_),
    .Y(_04185_));
 sky130_fd_sc_hd__o2bb2a_2 _18159_ (.A1_N(_04151_),
    .A2_N(_01973_),
    .B1(_04127_),
    .B2(_01978_),
    .X(_04186_));
 sky130_fd_sc_hd__o21ai_2 _18160_ (.A1(_04150_),
    .A2(_01972_),
    .B1(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__a31o_2 _18161_ (.A1(_04143_),
    .A2(_04184_),
    .A3(_04185_),
    .B1(_04187_),
    .X(_01979_));
 sky130_fd_sc_hd__or2_2 _18162_ (.A(_12889_),
    .B(_04179_),
    .X(_01980_));
 sky130_fd_sc_hd__buf_1 _18163_ (.A(_10617_),
    .X(_04188_));
 sky130_fd_sc_hd__or2_2 _18164_ (.A(_10886_),
    .B(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__o221a_2 _18165_ (.A1(_10854_),
    .A2(_04154_),
    .B1(_04139_),
    .B2(_11125_),
    .C1(_04189_),
    .X(_01984_));
 sky130_fd_sc_hd__a22o_2 _18166_ (.A1(_04103_),
    .A2(\timer[23] ),
    .B1(\irq_mask[23] ),
    .B2(_04104_),
    .X(_04190_));
 sky130_fd_sc_hd__a21oi_2 _18167_ (.A1(_04102_),
    .A2(\cpuregs_rs1[23] ),
    .B1(_04190_),
    .Y(_01986_));
 sky130_fd_sc_hd__o22a_2 _18168_ (.A1(_12556_),
    .A2(_12439_),
    .B1(\reg_pc[23] ),
    .B2(\decoded_imm[23] ),
    .X(_04191_));
 sky130_fd_sc_hd__o21ai_2 _18169_ (.A1(_12552_),
    .A2(_12438_),
    .B1(_04185_),
    .Y(_04192_));
 sky130_fd_sc_hd__nand2_2 _18170_ (.A(_04191_),
    .B(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__or2_2 _18171_ (.A(_04191_),
    .B(_04192_),
    .X(_04194_));
 sky130_fd_sc_hd__o2bb2a_2 _18172_ (.A1_N(_04151_),
    .A2_N(_01982_),
    .B1(_10470_),
    .B2(_01987_),
    .X(_04195_));
 sky130_fd_sc_hd__o21ai_2 _18173_ (.A1(_04150_),
    .A2(_01981_),
    .B1(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__a31o_2 _18174_ (.A1(_04143_),
    .A2(_04193_),
    .A3(_04194_),
    .B1(_04196_),
    .X(_01988_));
 sky130_fd_sc_hd__or2_2 _18175_ (.A(_12782_),
    .B(_04179_),
    .X(_01989_));
 sky130_fd_sc_hd__buf_1 _18176_ (.A(_10618_),
    .X(_04197_));
 sky130_fd_sc_hd__or2_2 _18177_ (.A(_10885_),
    .B(_04188_),
    .X(_04198_));
 sky130_fd_sc_hd__o221a_2 _18178_ (.A1(_10853_),
    .A2(_04154_),
    .B1(_04197_),
    .B2(_11124_),
    .C1(_04198_),
    .X(_01993_));
 sky130_fd_sc_hd__nand2_2 _18179_ (.A(_04141_),
    .B(\cpuregs_rs1[24] ),
    .Y(_04199_));
 sky130_fd_sc_hd__o221a_2 _18180_ (.A1(_11735_),
    .A2(_12427_),
    .B1(_10522_),
    .B2(_11741_),
    .C1(_04199_),
    .X(_01995_));
 sky130_fd_sc_hd__o21ai_2 _18181_ (.A1(_12556_),
    .A2(_12439_),
    .B1(_04193_),
    .Y(_04200_));
 sky130_fd_sc_hd__o22a_2 _18182_ (.A1(_12560_),
    .A2(_12440_),
    .B1(\reg_pc[24] ),
    .B2(\decoded_imm[24] ),
    .X(_04201_));
 sky130_fd_sc_hd__or2_2 _18183_ (.A(_04200_),
    .B(_04201_),
    .X(_04202_));
 sky130_fd_sc_hd__nand2_2 _18184_ (.A(_04200_),
    .B(_04201_),
    .Y(_04203_));
 sky130_fd_sc_hd__o2bb2a_2 _18185_ (.A1_N(_11084_),
    .A2_N(_01991_),
    .B1(_10470_),
    .B2(_01996_),
    .X(_04204_));
 sky130_fd_sc_hd__o21ai_2 _18186_ (.A1(_12781_),
    .A2(_01990_),
    .B1(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__a31o_2 _18187_ (.A1(_10604_),
    .A2(_04202_),
    .A3(_04203_),
    .B1(_04205_),
    .X(_01997_));
 sky130_fd_sc_hd__or2_2 _18188_ (.A(_12798_),
    .B(_04179_),
    .X(_01998_));
 sky130_fd_sc_hd__buf_1 _18189_ (.A(_10616_),
    .X(_04206_));
 sky130_fd_sc_hd__or2_2 _18190_ (.A(_10884_),
    .B(_04188_),
    .X(_04207_));
 sky130_fd_sc_hd__o221a_2 _18191_ (.A1(_10852_),
    .A2(_04206_),
    .B1(_04197_),
    .B2(_11123_),
    .C1(_04207_),
    .X(_02002_));
 sky130_fd_sc_hd__a22o_2 _18192_ (.A1(_12833_),
    .A2(\timer[25] ),
    .B1(\irq_mask[25] ),
    .B2(_12835_),
    .X(_04208_));
 sky130_fd_sc_hd__a21oi_2 _18193_ (.A1(_12804_),
    .A2(\cpuregs_rs1[25] ),
    .B1(_04208_),
    .Y(_02004_));
 sky130_fd_sc_hd__nor2_2 _18194_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .Y(_04209_));
 sky130_fd_sc_hd__a21oi_2 _18195_ (.A1(\reg_pc[25] ),
    .A2(\decoded_imm[25] ),
    .B1(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__o21ai_2 _18196_ (.A1(_12560_),
    .A2(_12440_),
    .B1(_04203_),
    .Y(_04211_));
 sky130_fd_sc_hd__or2_2 _18197_ (.A(_04210_),
    .B(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__a21oi_2 _18198_ (.A1(_04210_),
    .A2(_04211_),
    .B1(_12796_),
    .Y(_04213_));
 sky130_fd_sc_hd__o22ai_2 _18199_ (.A1(_12255_),
    .A2(_01999_),
    .B1(_12794_),
    .B2(_02005_),
    .Y(_04214_));
 sky130_fd_sc_hd__a221o_2 _18200_ (.A1(_12866_),
    .A2(_02000_),
    .B1(_04212_),
    .B2(_04213_),
    .C1(_04214_),
    .X(_02006_));
 sky130_fd_sc_hd__or2_2 _18201_ (.A(_12813_),
    .B(_04179_),
    .X(_02007_));
 sky130_fd_sc_hd__or2_2 _18202_ (.A(_10883_),
    .B(_04188_),
    .X(_04215_));
 sky130_fd_sc_hd__o221a_2 _18203_ (.A1(_10851_),
    .A2(_04206_),
    .B1(_04197_),
    .B2(_11122_),
    .C1(_04215_),
    .X(_02011_));
 sky130_fd_sc_hd__nand2_2 _18204_ (.A(_04141_),
    .B(\cpuregs_rs1[26] ),
    .Y(_04216_));
 sky130_fd_sc_hd__o221a_2 _18205_ (.A1(_11735_),
    .A2(_12377_),
    .B1(_10523_),
    .B2(_11741_),
    .C1(_04216_),
    .X(_02013_));
 sky130_fd_sc_hd__o32a_2 _18206_ (.A1(_12560_),
    .A2(_12440_),
    .A3(_04209_),
    .B1(_12564_),
    .B2(_12441_),
    .X(_04217_));
 sky130_vsdinv _18207_ (.A(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__a31o_2 _18208_ (.A1(_04201_),
    .A2(_04210_),
    .A3(_04200_),
    .B1(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__o22a_2 _18209_ (.A1(_12569_),
    .A2(_12442_),
    .B1(\reg_pc[26] ),
    .B2(\decoded_imm[26] ),
    .X(_04220_));
 sky130_fd_sc_hd__or2_2 _18210_ (.A(_04219_),
    .B(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__nand2_2 _18211_ (.A(_04219_),
    .B(_04220_),
    .Y(_04222_));
 sky130_fd_sc_hd__o2bb2a_2 _18212_ (.A1_N(_11084_),
    .A2_N(_02009_),
    .B1(_10470_),
    .B2(_02014_),
    .X(_04223_));
 sky130_fd_sc_hd__o21ai_2 _18213_ (.A1(_12781_),
    .A2(_02008_),
    .B1(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__a31o_2 _18214_ (.A1(_10604_),
    .A2(_04221_),
    .A3(_04222_),
    .B1(_04224_),
    .X(_02015_));
 sky130_fd_sc_hd__or2_2 _18215_ (.A(_12827_),
    .B(_04179_),
    .X(_02016_));
 sky130_fd_sc_hd__or2_2 _18216_ (.A(_10882_),
    .B(_04188_),
    .X(_04225_));
 sky130_fd_sc_hd__o221a_2 _18217_ (.A1(_10850_),
    .A2(_04206_),
    .B1(_04197_),
    .B2(_11121_),
    .C1(_04225_),
    .X(_02020_));
 sky130_fd_sc_hd__a22o_2 _18218_ (.A1(_12833_),
    .A2(\timer[27] ),
    .B1(\irq_mask[27] ),
    .B2(_12835_),
    .X(_04226_));
 sky130_fd_sc_hd__a21oi_2 _18219_ (.A1(_12804_),
    .A2(\cpuregs_rs1[27] ),
    .B1(_04226_),
    .Y(_02022_));
 sky130_fd_sc_hd__nor2_2 _18220_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .Y(_04227_));
 sky130_fd_sc_hd__a21oi_2 _18221_ (.A1(\reg_pc[27] ),
    .A2(\decoded_imm[27] ),
    .B1(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__o21ai_2 _18222_ (.A1(_12569_),
    .A2(_12442_),
    .B1(_04222_),
    .Y(_04229_));
 sky130_fd_sc_hd__or2_2 _18223_ (.A(_04228_),
    .B(_04229_),
    .X(_04230_));
 sky130_fd_sc_hd__a21oi_2 _18224_ (.A1(_04228_),
    .A2(_04229_),
    .B1(_12796_),
    .Y(_04231_));
 sky130_fd_sc_hd__o22ai_2 _18225_ (.A1(_12255_),
    .A2(_02017_),
    .B1(_12794_),
    .B2(_02023_),
    .Y(_04232_));
 sky130_fd_sc_hd__a221o_2 _18226_ (.A1(_12866_),
    .A2(_02018_),
    .B1(_04230_),
    .B2(_04231_),
    .C1(_04232_),
    .X(_02024_));
 sky130_fd_sc_hd__or2_2 _18227_ (.A(_12845_),
    .B(_12771_),
    .X(_02025_));
 sky130_fd_sc_hd__or2_2 _18228_ (.A(_10881_),
    .B(_04188_),
    .X(_04233_));
 sky130_fd_sc_hd__o221a_2 _18229_ (.A1(_10849_),
    .A2(_04206_),
    .B1(_04197_),
    .B2(_11120_),
    .C1(_04233_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_2 _18230_ (.A(_04141_),
    .B(\cpuregs_rs1[28] ),
    .Y(_04234_));
 sky130_fd_sc_hd__o221a_2 _18231_ (.A1(_11735_),
    .A2(_12429_),
    .B1(_10541_),
    .B2(_11741_),
    .C1(_04234_),
    .X(_02031_));
 sky130_fd_sc_hd__o2bb2a_2 _18232_ (.A1_N(_11085_),
    .A2_N(_02027_),
    .B1(_11031_),
    .B2(_02032_),
    .X(_04235_));
 sky130_fd_sc_hd__o32a_2 _18233_ (.A1(_12569_),
    .A2(_12442_),
    .A3(_04227_),
    .B1(_12576_),
    .B2(_12443_),
    .X(_04236_));
 sky130_vsdinv _18234_ (.A(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__a31o_2 _18235_ (.A1(_04220_),
    .A2(_04228_),
    .A3(_04219_),
    .B1(_04237_),
    .X(_04238_));
 sky130_fd_sc_hd__nor2_2 _18236_ (.A(\reg_pc[28] ),
    .B(\decoded_imm[28] ),
    .Y(_04239_));
 sky130_fd_sc_hd__a21oi_2 _18237_ (.A1(\reg_pc[28] ),
    .A2(\decoded_imm[28] ),
    .B1(_04239_),
    .Y(_04240_));
 sky130_vsdinv _18238_ (.A(_04238_),
    .Y(_04241_));
 sky130_vsdinv _18239_ (.A(_04240_),
    .Y(_04242_));
 sky130_fd_sc_hd__a221o_2 _18240_ (.A1(_04238_),
    .A2(_04240_),
    .B1(_04241_),
    .B2(_04242_),
    .C1(_10610_),
    .X(_04243_));
 sky130_fd_sc_hd__o211ai_2 _18241_ (.A1(_12256_),
    .A2(_02026_),
    .B1(_04235_),
    .C1(_04243_),
    .Y(_02033_));
 sky130_fd_sc_hd__or2_2 _18242_ (.A(_12857_),
    .B(_12771_),
    .X(_02034_));
 sky130_fd_sc_hd__or2_2 _18243_ (.A(_10880_),
    .B(_12861_),
    .X(_04244_));
 sky130_fd_sc_hd__o221a_2 _18244_ (.A1(_10848_),
    .A2(_04206_),
    .B1(_04197_),
    .B2(_11119_),
    .C1(_04244_),
    .X(_02038_));
 sky130_fd_sc_hd__a22o_2 _18245_ (.A1(_12833_),
    .A2(\timer[29] ),
    .B1(\irq_mask[29] ),
    .B2(_12835_),
    .X(_04245_));
 sky130_fd_sc_hd__a21oi_2 _18246_ (.A1(_12804_),
    .A2(\cpuregs_rs1[29] ),
    .B1(_04245_),
    .Y(_02040_));
 sky130_fd_sc_hd__o2bb2a_2 _18247_ (.A1_N(_11085_),
    .A2_N(_02036_),
    .B1(_11031_),
    .B2(_02041_),
    .X(_04246_));
 sky130_fd_sc_hd__o22a_2 _18248_ (.A1(_12580_),
    .A2(_12444_),
    .B1(_04241_),
    .B2(_04239_),
    .X(_04247_));
 sky130_vsdinv _18249_ (.A(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__nor2_2 _18250_ (.A(\reg_pc[29] ),
    .B(\decoded_imm[29] ),
    .Y(_04249_));
 sky130_fd_sc_hd__a21oi_2 _18251_ (.A1(\reg_pc[29] ),
    .A2(\decoded_imm[29] ),
    .B1(_04249_),
    .Y(_04250_));
 sky130_vsdinv _18252_ (.A(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__a221o_2 _18253_ (.A1(_04248_),
    .A2(_04250_),
    .B1(_04247_),
    .B2(_04251_),
    .C1(_10610_),
    .X(_04252_));
 sky130_fd_sc_hd__o211ai_2 _18254_ (.A1(_12809_),
    .A2(_02035_),
    .B1(_04246_),
    .C1(_04252_),
    .Y(_02042_));
 sky130_fd_sc_hd__or2_2 _18255_ (.A(_12873_),
    .B(_12771_),
    .X(_02043_));
 sky130_fd_sc_hd__or2_2 _18256_ (.A(_10879_),
    .B(_12861_),
    .X(_04253_));
 sky130_fd_sc_hd__o221a_2 _18257_ (.A1(_10847_),
    .A2(_04206_),
    .B1(_11773_),
    .B2(_11118_),
    .C1(_04253_),
    .X(_02047_));
 sky130_fd_sc_hd__nand2_2 _18258_ (.A(_12803_),
    .B(\cpuregs_rs1[30] ),
    .Y(_04254_));
 sky130_fd_sc_hd__o221a_2 _18259_ (.A1(_11735_),
    .A2(_12431_),
    .B1(_10542_),
    .B2(_11741_),
    .C1(_04254_),
    .X(_02049_));
 sky130_fd_sc_hd__o22a_2 _18260_ (.A1(_12594_),
    .A2(_12446_),
    .B1(\reg_pc[30] ),
    .B2(\decoded_imm[30] ),
    .X(_04255_));
 sky130_fd_sc_hd__o22ai_2 _18261_ (.A1(_12589_),
    .A2(_12445_),
    .B1(_04247_),
    .B2(_04249_),
    .Y(_04256_));
 sky130_fd_sc_hd__or2_2 _18262_ (.A(_04255_),
    .B(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__nand2_2 _18263_ (.A(_04255_),
    .B(_04256_),
    .Y(_04258_));
 sky130_fd_sc_hd__o2bb2a_2 _18264_ (.A1_N(_11084_),
    .A2_N(_02045_),
    .B1(_10470_),
    .B2(_02050_),
    .X(_04259_));
 sky130_fd_sc_hd__o21ai_2 _18265_ (.A1(_12781_),
    .A2(_02044_),
    .B1(_04259_),
    .Y(_04260_));
 sky130_fd_sc_hd__a31o_2 _18266_ (.A1(_10604_),
    .A2(_04257_),
    .A3(_04258_),
    .B1(_04260_),
    .X(_02051_));
 sky130_fd_sc_hd__or2_2 _18267_ (.A(_12888_),
    .B(_12771_),
    .X(_02052_));
 sky130_fd_sc_hd__or2_2 _18268_ (.A(_10878_),
    .B(_12861_),
    .X(_04261_));
 sky130_fd_sc_hd__o221a_2 _18269_ (.A1(_10973_),
    .A2(_11766_),
    .B1(_11773_),
    .B2(_11210_),
    .C1(_04261_),
    .X(_02056_));
 sky130_fd_sc_hd__a22o_2 _18270_ (.A1(_12833_),
    .A2(\timer[31] ),
    .B1(\irq_mask[31] ),
    .B2(_12835_),
    .X(_04262_));
 sky130_fd_sc_hd__a21oi_2 _18271_ (.A1(_12804_),
    .A2(\cpuregs_rs1[31] ),
    .B1(_04262_),
    .Y(_02058_));
 sky130_fd_sc_hd__o21ai_2 _18272_ (.A1(_12594_),
    .A2(_12446_),
    .B1(_04258_),
    .Y(_04263_));
 sky130_fd_sc_hd__a221o_2 _18273_ (.A1(\reg_pc[31] ),
    .A2(_12173_),
    .B1(_12599_),
    .B2(\decoded_imm[31] ),
    .C1(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__o221ai_2 _18274_ (.A1(\reg_pc[31] ),
    .A2(\decoded_imm[31] ),
    .B1(_12599_),
    .B2(_12173_),
    .C1(_04263_),
    .Y(_04265_));
 sky130_fd_sc_hd__o2bb2a_2 _18275_ (.A1_N(_11084_),
    .A2_N(_02054_),
    .B1(_10470_),
    .B2(_02059_),
    .X(_04266_));
 sky130_fd_sc_hd__o21ai_2 _18276_ (.A1(_12781_),
    .A2(_02053_),
    .B1(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__a31o_2 _18277_ (.A1(_10604_),
    .A2(_04264_),
    .A3(_04265_),
    .B1(_04267_),
    .X(_02060_));
 sky130_fd_sc_hd__or2_2 _18278_ (.A(\decoded_rd[4] ),
    .B(_00308_),
    .X(_02061_));
 sky130_vsdinv _18279_ (.A(_12211_),
    .Y(_02062_));
 sky130_fd_sc_hd__o21ai_2 _18280_ (.A1(_12274_),
    .A2(_02064_),
    .B1(_12369_),
    .Y(_02065_));
 sky130_fd_sc_hd__nor3_2 _18281_ (.A(_10564_),
    .B(_02410_),
    .C(_00308_),
    .Y(_02066_));
 sky130_fd_sc_hd__buf_1 _18282_ (.A(_01706_),
    .X(_02067_));
 sky130_fd_sc_hd__nor2_2 _18283_ (.A(_10786_),
    .B(_12368_),
    .Y(_04268_));
 sky130_fd_sc_hd__o211ai_2 _18284_ (.A1(_12274_),
    .A2(_04268_),
    .B1(_12369_),
    .C1(_12256_),
    .Y(_02068_));
 sky130_fd_sc_hd__buf_1 _18285_ (.A(_10649_),
    .X(_04269_));
 sky130_fd_sc_hd__or2_2 _18286_ (.A(latched_branch),
    .B(_11256_),
    .X(_04270_));
 sky130_fd_sc_hd__and3_2 _18287_ (.A(_04269_),
    .B(_10648_),
    .C(_04270_),
    .X(_02069_));
 sky130_vsdinv _18288_ (.A(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__buf_1 _18289_ (.A(_04271_),
    .X(_04272_));
 sky130_fd_sc_hd__a22o_2 _18290_ (.A1(_02070_),
    .A2(_04272_),
    .B1(_10655_),
    .B2(\reg_next_pc[0] ),
    .X(_04273_));
 sky130_fd_sc_hd__a31o_2 _18291_ (.A1(_11079_),
    .A2(\irq_pending[0] ),
    .A3(_10645_),
    .B1(_04273_),
    .X(_02071_));
 sky130_fd_sc_hd__buf_1 _18292_ (.A(_04272_),
    .X(_04274_));
 sky130_fd_sc_hd__and3_2 _18293_ (.A(_10510_),
    .B(\irq_pending[1] ),
    .C(_10645_),
    .X(_04275_));
 sky130_fd_sc_hd__a221o_2 _18294_ (.A1(_01465_),
    .A2(_04274_),
    .B1(_10656_),
    .B2(\reg_next_pc[1] ),
    .C1(_04275_),
    .X(_02072_));
 sky130_fd_sc_hd__and3_2 _18295_ (.A(_10511_),
    .B(\irq_pending[2] ),
    .C(_10645_),
    .X(_04276_));
 sky130_fd_sc_hd__a221o_2 _18296_ (.A1(_00293_),
    .A2(_04274_),
    .B1(_10656_),
    .B2(\reg_next_pc[2] ),
    .C1(_04276_),
    .X(_02074_));
 sky130_fd_sc_hd__nor2_2 _18297_ (.A(_12458_),
    .B(_02073_),
    .Y(_04277_));
 sky130_fd_sc_hd__a21oi_2 _18298_ (.A1(_12458_),
    .A2(_02073_),
    .B1(_04277_),
    .Y(_02075_));
 sky130_fd_sc_hd__nor3_2 _18299_ (.A(\irq_mask[3] ),
    .B(_10513_),
    .C(_04269_),
    .Y(_04278_));
 sky130_fd_sc_hd__a221o_2 _18300_ (.A1(_01468_),
    .A2(_04274_),
    .B1(_10656_),
    .B2(\reg_next_pc[3] ),
    .C1(_04278_),
    .X(_02076_));
 sky130_fd_sc_hd__nand2_2 _18301_ (.A(\reg_pc[4] ),
    .B(_04277_),
    .Y(_04279_));
 sky130_fd_sc_hd__o21a_2 _18302_ (.A1(\reg_pc[4] ),
    .A2(_04277_),
    .B1(_04279_),
    .X(_02077_));
 sky130_fd_sc_hd__nor3_2 _18303_ (.A(\irq_mask[4] ),
    .B(_10530_),
    .C(_04269_),
    .Y(_04280_));
 sky130_fd_sc_hd__a221o_2 _18304_ (.A1(_01472_),
    .A2(_04274_),
    .B1(_10656_),
    .B2(\reg_next_pc[4] ),
    .C1(_04280_),
    .X(_02078_));
 sky130_fd_sc_hd__nor2_2 _18305_ (.A(_12468_),
    .B(_04279_),
    .Y(_04281_));
 sky130_fd_sc_hd__a21oi_2 _18306_ (.A1(_12468_),
    .A2(_04279_),
    .B1(_04281_),
    .Y(_02079_));
 sky130_fd_sc_hd__buf_1 _18307_ (.A(_10654_),
    .X(_04282_));
 sky130_fd_sc_hd__and3_2 _18308_ (.A(_10528_),
    .B(\irq_pending[5] ),
    .C(_10645_),
    .X(_04283_));
 sky130_fd_sc_hd__a221o_2 _18309_ (.A1(_01476_),
    .A2(_04274_),
    .B1(_04282_),
    .B2(\reg_next_pc[5] ),
    .C1(_04283_),
    .X(_02080_));
 sky130_fd_sc_hd__nand2_2 _18310_ (.A(\reg_pc[6] ),
    .B(_04281_),
    .Y(_04284_));
 sky130_fd_sc_hd__o21a_2 _18311_ (.A1(\reg_pc[6] ),
    .A2(_04281_),
    .B1(_04284_),
    .X(_02081_));
 sky130_fd_sc_hd__nor3_2 _18312_ (.A(\irq_mask[6] ),
    .B(_10531_),
    .C(_04269_),
    .Y(_04285_));
 sky130_fd_sc_hd__a221o_2 _18313_ (.A1(_01479_),
    .A2(_04274_),
    .B1(_04282_),
    .B2(\reg_next_pc[6] ),
    .C1(_04285_),
    .X(_02082_));
 sky130_fd_sc_hd__or2_2 _18314_ (.A(_12478_),
    .B(_04284_),
    .X(_04286_));
 sky130_vsdinv _18315_ (.A(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__a21oi_2 _18316_ (.A1(_12478_),
    .A2(_04284_),
    .B1(_04287_),
    .Y(_02083_));
 sky130_fd_sc_hd__buf_1 _18317_ (.A(_04272_),
    .X(_04288_));
 sky130_fd_sc_hd__and3_2 _18318_ (.A(_10529_),
    .B(\irq_pending[7] ),
    .C(_10645_),
    .X(_04289_));
 sky130_fd_sc_hd__a221o_2 _18319_ (.A1(_01482_),
    .A2(_04288_),
    .B1(_04282_),
    .B2(\reg_next_pc[7] ),
    .C1(_04289_),
    .X(_02084_));
 sky130_fd_sc_hd__or2_2 _18320_ (.A(_12483_),
    .B(_04286_),
    .X(_04290_));
 sky130_fd_sc_hd__o21a_2 _18321_ (.A1(\reg_pc[8] ),
    .A2(_04287_),
    .B1(_04290_),
    .X(_02085_));
 sky130_fd_sc_hd__nor3_2 _18322_ (.A(\irq_mask[8] ),
    .B(_10549_),
    .C(_04269_),
    .Y(_04291_));
 sky130_fd_sc_hd__a221o_2 _18323_ (.A1(_01485_),
    .A2(_04288_),
    .B1(_04282_),
    .B2(\reg_next_pc[8] ),
    .C1(_04291_),
    .X(_02086_));
 sky130_fd_sc_hd__or2_2 _18324_ (.A(_12492_),
    .B(_04290_),
    .X(_04292_));
 sky130_vsdinv _18325_ (.A(_04292_),
    .Y(_04293_));
 sky130_fd_sc_hd__a21oi_2 _18326_ (.A1(_12492_),
    .A2(_04290_),
    .B1(_04293_),
    .Y(_02087_));
 sky130_fd_sc_hd__buf_1 _18327_ (.A(\irq_state[1] ),
    .X(_04294_));
 sky130_fd_sc_hd__buf_1 _18328_ (.A(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__and3_2 _18329_ (.A(_10547_),
    .B(\irq_pending[9] ),
    .C(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__a221o_2 _18330_ (.A1(_01488_),
    .A2(_04288_),
    .B1(_04282_),
    .B2(\reg_next_pc[9] ),
    .C1(_04296_),
    .X(_02088_));
 sky130_fd_sc_hd__or2_2 _18331_ (.A(_12496_),
    .B(_04292_),
    .X(_04297_));
 sky130_fd_sc_hd__o21a_2 _18332_ (.A1(\reg_pc[10] ),
    .A2(_04293_),
    .B1(_04297_),
    .X(_02089_));
 sky130_fd_sc_hd__nor3_2 _18333_ (.A(\irq_mask[10] ),
    .B(_10550_),
    .C(_04269_),
    .Y(_04298_));
 sky130_fd_sc_hd__a221o_2 _18334_ (.A1(_01491_),
    .A2(_04288_),
    .B1(_04282_),
    .B2(\reg_next_pc[10] ),
    .C1(_04298_),
    .X(_02090_));
 sky130_fd_sc_hd__or2_2 _18335_ (.A(_12502_),
    .B(_04297_),
    .X(_04299_));
 sky130_vsdinv _18336_ (.A(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__a21oi_2 _18337_ (.A1(_12502_),
    .A2(_04297_),
    .B1(_04300_),
    .Y(_02091_));
 sky130_fd_sc_hd__buf_1 _18338_ (.A(_10654_),
    .X(_04301_));
 sky130_fd_sc_hd__and3_2 _18339_ (.A(_10548_),
    .B(\irq_pending[11] ),
    .C(_04295_),
    .X(_04302_));
 sky130_fd_sc_hd__a221o_2 _18340_ (.A1(_01494_),
    .A2(_04288_),
    .B1(_04301_),
    .B2(\reg_next_pc[11] ),
    .C1(_04302_),
    .X(_02092_));
 sky130_fd_sc_hd__or2_2 _18341_ (.A(_12506_),
    .B(_04299_),
    .X(_04303_));
 sky130_fd_sc_hd__o21a_2 _18342_ (.A1(\reg_pc[12] ),
    .A2(_04300_),
    .B1(_04303_),
    .X(_02093_));
 sky130_fd_sc_hd__buf_1 _18343_ (.A(_10649_),
    .X(_04304_));
 sky130_fd_sc_hd__nor3_2 _18344_ (.A(\irq_mask[12] ),
    .B(_10537_),
    .C(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__a221o_2 _18345_ (.A1(_01497_),
    .A2(_04288_),
    .B1(_04301_),
    .B2(\reg_next_pc[12] ),
    .C1(_04305_),
    .X(_02094_));
 sky130_fd_sc_hd__or2_2 _18346_ (.A(_12510_),
    .B(_04303_),
    .X(_04306_));
 sky130_vsdinv _18347_ (.A(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__a21oi_2 _18348_ (.A1(_12510_),
    .A2(_04303_),
    .B1(_04307_),
    .Y(_02095_));
 sky130_fd_sc_hd__buf_1 _18349_ (.A(_04272_),
    .X(_04308_));
 sky130_fd_sc_hd__and3_2 _18350_ (.A(_10535_),
    .B(\irq_pending[13] ),
    .C(_04295_),
    .X(_04309_));
 sky130_fd_sc_hd__a221o_2 _18351_ (.A1(_01500_),
    .A2(_04308_),
    .B1(_04301_),
    .B2(\reg_next_pc[13] ),
    .C1(_04309_),
    .X(_02096_));
 sky130_fd_sc_hd__or2_2 _18352_ (.A(_12515_),
    .B(_04306_),
    .X(_04310_));
 sky130_fd_sc_hd__o21a_2 _18353_ (.A1(\reg_pc[14] ),
    .A2(_04307_),
    .B1(_04310_),
    .X(_02097_));
 sky130_fd_sc_hd__nor3_2 _18354_ (.A(\irq_mask[14] ),
    .B(_10538_),
    .C(_04304_),
    .Y(_04311_));
 sky130_fd_sc_hd__a221o_2 _18355_ (.A1(_01503_),
    .A2(_04308_),
    .B1(_04301_),
    .B2(\reg_next_pc[14] ),
    .C1(_04311_),
    .X(_02098_));
 sky130_fd_sc_hd__or2_2 _18356_ (.A(_12519_),
    .B(_04310_),
    .X(_04312_));
 sky130_vsdinv _18357_ (.A(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__a21oi_2 _18358_ (.A1(_12519_),
    .A2(_04310_),
    .B1(_04313_),
    .Y(_02099_));
 sky130_fd_sc_hd__and3_2 _18359_ (.A(_10536_),
    .B(\irq_pending[15] ),
    .C(_04295_),
    .X(_04314_));
 sky130_fd_sc_hd__a221o_2 _18360_ (.A1(_01506_),
    .A2(_04308_),
    .B1(_04301_),
    .B2(\reg_next_pc[15] ),
    .C1(_04314_),
    .X(_02100_));
 sky130_fd_sc_hd__or2_2 _18361_ (.A(_12523_),
    .B(_04312_),
    .X(_04315_));
 sky130_fd_sc_hd__o21a_2 _18362_ (.A1(\reg_pc[16] ),
    .A2(_04313_),
    .B1(_04315_),
    .X(_02101_));
 sky130_fd_sc_hd__nor3_2 _18363_ (.A(\irq_mask[16] ),
    .B(_10518_),
    .C(_04304_),
    .Y(_04316_));
 sky130_fd_sc_hd__a221o_2 _18364_ (.A1(_01509_),
    .A2(_04308_),
    .B1(_04301_),
    .B2(\reg_next_pc[16] ),
    .C1(_04316_),
    .X(_02102_));
 sky130_fd_sc_hd__or2_2 _18365_ (.A(_12529_),
    .B(_04315_),
    .X(_04317_));
 sky130_vsdinv _18366_ (.A(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__a21oi_2 _18367_ (.A1(_12529_),
    .A2(_04315_),
    .B1(_04318_),
    .Y(_02103_));
 sky130_fd_sc_hd__buf_1 _18368_ (.A(_10654_),
    .X(_04319_));
 sky130_fd_sc_hd__nor3_2 _18369_ (.A(\irq_mask[17] ),
    .B(_10516_),
    .C(_04304_),
    .Y(_04320_));
 sky130_fd_sc_hd__a221o_2 _18370_ (.A1(_01512_),
    .A2(_04308_),
    .B1(_04319_),
    .B2(\reg_next_pc[17] ),
    .C1(_04320_),
    .X(_02104_));
 sky130_fd_sc_hd__or2_2 _18371_ (.A(_12533_),
    .B(_04317_),
    .X(_04321_));
 sky130_fd_sc_hd__o21a_2 _18372_ (.A1(\reg_pc[18] ),
    .A2(_04318_),
    .B1(_04321_),
    .X(_02105_));
 sky130_fd_sc_hd__and3_2 _18373_ (.A(_11052_),
    .B(\irq_pending[18] ),
    .C(_04295_),
    .X(_04322_));
 sky130_fd_sc_hd__a221o_2 _18374_ (.A1(_01515_),
    .A2(_04308_),
    .B1(_04319_),
    .B2(\reg_next_pc[18] ),
    .C1(_04322_),
    .X(_02106_));
 sky130_fd_sc_hd__or2_2 _18375_ (.A(_12539_),
    .B(_04321_),
    .X(_04323_));
 sky130_vsdinv _18376_ (.A(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__a21oi_2 _18377_ (.A1(_12539_),
    .A2(_04321_),
    .B1(_04324_),
    .Y(_02107_));
 sky130_fd_sc_hd__buf_1 _18378_ (.A(_04272_),
    .X(_04325_));
 sky130_fd_sc_hd__nor3_2 _18379_ (.A(\irq_mask[19] ),
    .B(_10517_),
    .C(_04304_),
    .Y(_04326_));
 sky130_fd_sc_hd__a221o_2 _18380_ (.A1(_01518_),
    .A2(_04325_),
    .B1(_04319_),
    .B2(\reg_next_pc[19] ),
    .C1(_04326_),
    .X(_02108_));
 sky130_fd_sc_hd__or2_2 _18381_ (.A(_12544_),
    .B(_04323_),
    .X(_04327_));
 sky130_fd_sc_hd__o21a_2 _18382_ (.A1(\reg_pc[20] ),
    .A2(_04324_),
    .B1(_04327_),
    .X(_02109_));
 sky130_fd_sc_hd__and3_2 _18383_ (.A(_10553_),
    .B(\irq_pending[20] ),
    .C(_04295_),
    .X(_04328_));
 sky130_fd_sc_hd__a221o_2 _18384_ (.A1(_01521_),
    .A2(_04325_),
    .B1(_04319_),
    .B2(\reg_next_pc[20] ),
    .C1(_04328_),
    .X(_02110_));
 sky130_fd_sc_hd__or2_2 _18385_ (.A(_12548_),
    .B(_04327_),
    .X(_04329_));
 sky130_vsdinv _18386_ (.A(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__a21oi_2 _18387_ (.A1(_12548_),
    .A2(_04327_),
    .B1(_04330_),
    .Y(_02111_));
 sky130_fd_sc_hd__nor3_2 _18388_ (.A(\irq_mask[21] ),
    .B(_10555_),
    .C(_04304_),
    .Y(_04331_));
 sky130_fd_sc_hd__a221o_2 _18389_ (.A1(_01524_),
    .A2(_04325_),
    .B1(_04319_),
    .B2(\reg_next_pc[21] ),
    .C1(_04331_),
    .X(_02112_));
 sky130_fd_sc_hd__or2_2 _18390_ (.A(_12552_),
    .B(_04329_),
    .X(_04332_));
 sky130_fd_sc_hd__o21a_2 _18391_ (.A1(\reg_pc[22] ),
    .A2(_04330_),
    .B1(_04332_),
    .X(_02113_));
 sky130_fd_sc_hd__and3_2 _18392_ (.A(_10554_),
    .B(\irq_pending[22] ),
    .C(_04294_),
    .X(_04333_));
 sky130_fd_sc_hd__a221o_2 _18393_ (.A1(_01527_),
    .A2(_04325_),
    .B1(_04319_),
    .B2(\reg_next_pc[22] ),
    .C1(_04333_),
    .X(_02114_));
 sky130_fd_sc_hd__or2_2 _18394_ (.A(_12556_),
    .B(_04332_),
    .X(_04334_));
 sky130_vsdinv _18395_ (.A(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__a21oi_2 _18396_ (.A1(_12556_),
    .A2(_04332_),
    .B1(_04335_),
    .Y(_02115_));
 sky130_fd_sc_hd__buf_1 _18397_ (.A(_10654_),
    .X(_04336_));
 sky130_fd_sc_hd__nor3_2 _18398_ (.A(\irq_mask[23] ),
    .B(_10556_),
    .C(_10650_),
    .Y(_04337_));
 sky130_fd_sc_hd__a221o_2 _18399_ (.A1(_01530_),
    .A2(_04325_),
    .B1(_04336_),
    .B2(\reg_next_pc[23] ),
    .C1(_04337_),
    .X(_02116_));
 sky130_fd_sc_hd__or2_2 _18400_ (.A(_12560_),
    .B(_04334_),
    .X(_04338_));
 sky130_fd_sc_hd__o21a_2 _18401_ (.A1(\reg_pc[24] ),
    .A2(_04335_),
    .B1(_04338_),
    .X(_02117_));
 sky130_fd_sc_hd__and3_2 _18402_ (.A(_10522_),
    .B(\irq_pending[24] ),
    .C(_04294_),
    .X(_04339_));
 sky130_fd_sc_hd__a221o_2 _18403_ (.A1(_01533_),
    .A2(_04325_),
    .B1(_04336_),
    .B2(\reg_next_pc[24] ),
    .C1(_04339_),
    .X(_02118_));
 sky130_fd_sc_hd__or2_2 _18404_ (.A(_12564_),
    .B(_04338_),
    .X(_04340_));
 sky130_vsdinv _18405_ (.A(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__a21oi_2 _18406_ (.A1(_12564_),
    .A2(_04338_),
    .B1(_04341_),
    .Y(_02119_));
 sky130_fd_sc_hd__buf_1 _18407_ (.A(_04271_),
    .X(_04342_));
 sky130_fd_sc_hd__nor3_2 _18408_ (.A(\irq_mask[25] ),
    .B(_10524_),
    .C(_10650_),
    .Y(_04343_));
 sky130_fd_sc_hd__a221o_2 _18409_ (.A1(_01536_),
    .A2(_04342_),
    .B1(_04336_),
    .B2(\reg_next_pc[25] ),
    .C1(_04343_),
    .X(_02120_));
 sky130_fd_sc_hd__or2_2 _18410_ (.A(_12569_),
    .B(_04340_),
    .X(_04344_));
 sky130_fd_sc_hd__o21a_2 _18411_ (.A1(\reg_pc[26] ),
    .A2(_04341_),
    .B1(_04344_),
    .X(_02121_));
 sky130_fd_sc_hd__and3_2 _18412_ (.A(_10523_),
    .B(\irq_pending[26] ),
    .C(_04294_),
    .X(_04345_));
 sky130_fd_sc_hd__a221o_2 _18413_ (.A1(_01539_),
    .A2(_04342_),
    .B1(_04336_),
    .B2(\reg_next_pc[26] ),
    .C1(_04345_),
    .X(_02122_));
 sky130_fd_sc_hd__or2_2 _18414_ (.A(_12576_),
    .B(_04344_),
    .X(_04346_));
 sky130_vsdinv _18415_ (.A(_04346_),
    .Y(_04347_));
 sky130_fd_sc_hd__a21oi_2 _18416_ (.A1(_12576_),
    .A2(_04344_),
    .B1(_04347_),
    .Y(_02123_));
 sky130_fd_sc_hd__nor3_2 _18417_ (.A(\irq_mask[27] ),
    .B(_10525_),
    .C(_10650_),
    .Y(_04348_));
 sky130_fd_sc_hd__a221o_2 _18418_ (.A1(_01542_),
    .A2(_04342_),
    .B1(_04336_),
    .B2(\reg_next_pc[27] ),
    .C1(_04348_),
    .X(_02124_));
 sky130_fd_sc_hd__or2_2 _18419_ (.A(_12580_),
    .B(_04346_),
    .X(_04349_));
 sky130_fd_sc_hd__o21a_2 _18420_ (.A1(\reg_pc[28] ),
    .A2(_04347_),
    .B1(_04349_),
    .X(_02125_));
 sky130_fd_sc_hd__and3_2 _18421_ (.A(_10541_),
    .B(\irq_pending[28] ),
    .C(_04294_),
    .X(_04350_));
 sky130_fd_sc_hd__a221o_2 _18422_ (.A1(_01545_),
    .A2(_04342_),
    .B1(_04336_),
    .B2(\reg_next_pc[28] ),
    .C1(_04350_),
    .X(_02126_));
 sky130_fd_sc_hd__or2_2 _18423_ (.A(_12589_),
    .B(_04349_),
    .X(_04351_));
 sky130_vsdinv _18424_ (.A(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__a21oi_2 _18425_ (.A1(_12589_),
    .A2(_04349_),
    .B1(_04352_),
    .Y(_02127_));
 sky130_fd_sc_hd__nor3_2 _18426_ (.A(\irq_mask[29] ),
    .B(_10543_),
    .C(_10650_),
    .Y(_04353_));
 sky130_fd_sc_hd__a221o_2 _18427_ (.A1(_01548_),
    .A2(_04342_),
    .B1(_10655_),
    .B2(\reg_next_pc[29] ),
    .C1(_04353_),
    .X(_02128_));
 sky130_fd_sc_hd__or2_2 _18428_ (.A(_12594_),
    .B(_04351_),
    .X(_04354_));
 sky130_fd_sc_hd__o21a_2 _18429_ (.A1(\reg_pc[30] ),
    .A2(_04352_),
    .B1(_04354_),
    .X(_02129_));
 sky130_fd_sc_hd__and3_2 _18430_ (.A(_10542_),
    .B(\irq_pending[30] ),
    .C(_04294_),
    .X(_04355_));
 sky130_fd_sc_hd__a221o_2 _18431_ (.A1(_01551_),
    .A2(_04342_),
    .B1(_10655_),
    .B2(\reg_next_pc[30] ),
    .C1(_04355_),
    .X(_02130_));
 sky130_fd_sc_hd__a32o_2 _18432_ (.A1(\reg_pc[30] ),
    .A2(_04352_),
    .A3(_12599_),
    .B1(\reg_pc[31] ),
    .B2(_04354_),
    .X(_02131_));
 sky130_fd_sc_hd__nor3_2 _18433_ (.A(\irq_mask[31] ),
    .B(_10544_),
    .C(_10650_),
    .Y(_04356_));
 sky130_fd_sc_hd__a221o_2 _18434_ (.A1(_01554_),
    .A2(_04272_),
    .B1(_10655_),
    .B2(\reg_next_pc[31] ),
    .C1(_04356_),
    .X(_02132_));
 sky130_fd_sc_hd__or2_2 _18435_ (.A(instr_xor),
    .B(instr_xori),
    .X(_04357_));
 sky130_fd_sc_hd__buf_1 _18436_ (.A(_04357_),
    .X(_04358_));
 sky130_fd_sc_hd__or3_2 _18437_ (.A(is_compare),
    .B(_04358_),
    .C(_10631_),
    .X(_04359_));
 sky130_fd_sc_hd__nor2_2 _18438_ (.A(instr_and),
    .B(instr_andi),
    .Y(_04360_));
 sky130_fd_sc_hd__buf_1 _18439_ (.A(_04360_),
    .X(_04361_));
 sky130_fd_sc_hd__buf_1 _18440_ (.A(_04361_),
    .X(_04362_));
 sky130_fd_sc_hd__nor2_2 _18441_ (.A(instr_or),
    .B(instr_ori),
    .Y(_04363_));
 sky130_fd_sc_hd__buf_1 _18442_ (.A(_04363_),
    .X(_04364_));
 sky130_fd_sc_hd__buf_1 _18443_ (.A(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__or2_2 _18444_ (.A(instr_sll),
    .B(instr_slli),
    .X(_04366_));
 sky130_vsdinv _18445_ (.A(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__and4b_2 _18446_ (.A_N(_04359_),
    .B(_04362_),
    .C(_04365_),
    .D(_04367_),
    .X(_02133_));
 sky130_fd_sc_hd__buf_1 _18447_ (.A(_04357_),
    .X(_04368_));
 sky130_fd_sc_hd__buf_1 _18448_ (.A(_10631_),
    .X(_04369_));
 sky130_vsdinv _18449_ (.A(is_compare),
    .Y(_04370_));
 sky130_fd_sc_hd__nor2_2 _18450_ (.A(_11364_),
    .B(_11863_),
    .Y(_04371_));
 sky130_vsdinv _18451_ (.A(\alu_shl[0] ),
    .Y(_04372_));
 sky130_fd_sc_hd__o32a_2 _18452_ (.A1(_12281_),
    .A2(_12196_),
    .A3(_04361_),
    .B1(_04372_),
    .B2(_04367_),
    .X(_04373_));
 sky130_fd_sc_hd__o221ai_2 _18453_ (.A1(_00343_),
    .A2(_04370_),
    .B1(_04365_),
    .B2(_04371_),
    .C1(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__a221o_2 _18454_ (.A1(_02591_),
    .A2(_04368_),
    .B1(\alu_shr[0] ),
    .B2(_04369_),
    .C1(_04374_),
    .X(_02134_));
 sky130_fd_sc_hd__buf_1 _18455_ (.A(_04369_),
    .X(_04375_));
 sky130_fd_sc_hd__buf_1 _18456_ (.A(_04366_),
    .X(_04376_));
 sky130_fd_sc_hd__buf_1 _18457_ (.A(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__a22o_2 _18458_ (.A1(\alu_shl[1] ),
    .A2(_04377_),
    .B1(_12325_),
    .B2(_04368_),
    .X(_04378_));
 sky130_fd_sc_hd__o32a_2 _18459_ (.A1(_02318_),
    .A2(_12770_),
    .A3(_04362_),
    .B1(_12324_),
    .B2(_04365_),
    .X(_04379_));
 sky130_vsdinv _18460_ (.A(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__a211o_2 _18461_ (.A1(\alu_shr[1] ),
    .A2(_04375_),
    .B1(_04378_),
    .C1(_04380_),
    .X(_02135_));
 sky130_fd_sc_hd__a22o_2 _18462_ (.A1(\alu_shl[2] ),
    .A2(_04377_),
    .B1(_12334_),
    .B2(_04368_),
    .X(_04381_));
 sky130_fd_sc_hd__o32a_2 _18463_ (.A1(_12191_),
    .A2(_12459_),
    .A3(_04362_),
    .B1(_12333_),
    .B2(_04365_),
    .X(_04382_));
 sky130_vsdinv _18464_ (.A(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__a211o_2 _18465_ (.A1(\alu_shr[2] ),
    .A2(_04375_),
    .B1(_04381_),
    .C1(_04383_),
    .X(_02136_));
 sky130_fd_sc_hd__a22o_2 _18466_ (.A1(\alu_shl[3] ),
    .A2(_04377_),
    .B1(_12327_),
    .B2(_04368_),
    .X(_04384_));
 sky130_fd_sc_hd__o32a_2 _18467_ (.A1(_12187_),
    .A2(_12464_),
    .A3(_04362_),
    .B1(_12326_),
    .B2(_04365_),
    .X(_04385_));
 sky130_vsdinv _18468_ (.A(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__a211o_2 _18469_ (.A1(\alu_shr[3] ),
    .A2(_04375_),
    .B1(_04384_),
    .C1(_04386_),
    .X(_02137_));
 sky130_fd_sc_hd__a22o_2 _18470_ (.A1(\alu_shl[4] ),
    .A2(_04377_),
    .B1(_12330_),
    .B2(_04368_),
    .X(_04387_));
 sky130_fd_sc_hd__o32a_2 _18471_ (.A1(_12185_),
    .A2(_12469_),
    .A3(_04362_),
    .B1(_12329_),
    .B2(_04365_),
    .X(_04388_));
 sky130_vsdinv _18472_ (.A(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__a211o_2 _18473_ (.A1(\alu_shr[4] ),
    .A2(_04375_),
    .B1(_04387_),
    .C1(_04389_),
    .X(_02138_));
 sky130_fd_sc_hd__a22o_2 _18474_ (.A1(\alu_shl[5] ),
    .A2(_04377_),
    .B1(_12321_),
    .B2(_04368_),
    .X(_04390_));
 sky130_fd_sc_hd__inv_2 _18475_ (.A(mem_la_wdata[5]),
    .Y(_02330_));
 sky130_fd_sc_hd__buf_1 _18476_ (.A(_04364_),
    .X(_04391_));
 sky130_fd_sc_hd__o32a_2 _18477_ (.A1(_02330_),
    .A2(_12474_),
    .A3(_04362_),
    .B1(_12320_),
    .B2(_04391_),
    .X(_04392_));
 sky130_vsdinv _18478_ (.A(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__a211o_2 _18479_ (.A1(\alu_shr[5] ),
    .A2(_04375_),
    .B1(_04390_),
    .C1(_04393_),
    .X(_02139_));
 sky130_fd_sc_hd__buf_1 _18480_ (.A(_04358_),
    .X(_04394_));
 sky130_fd_sc_hd__a22o_2 _18481_ (.A1(\alu_shl[6] ),
    .A2(_04377_),
    .B1(_12332_),
    .B2(_04394_),
    .X(_04395_));
 sky130_fd_sc_hd__inv_2 _18482_ (.A(_11358_),
    .Y(_02333_));
 sky130_fd_sc_hd__buf_1 _18483_ (.A(_04361_),
    .X(_04396_));
 sky130_fd_sc_hd__o32a_2 _18484_ (.A1(_02333_),
    .A2(_12476_),
    .A3(_04396_),
    .B1(_12331_),
    .B2(_04391_),
    .X(_04397_));
 sky130_vsdinv _18485_ (.A(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__a211o_2 _18486_ (.A1(\alu_shr[6] ),
    .A2(_04375_),
    .B1(_04395_),
    .C1(_04398_),
    .X(_02140_));
 sky130_fd_sc_hd__buf_1 _18487_ (.A(_04369_),
    .X(_04399_));
 sky130_fd_sc_hd__buf_1 _18488_ (.A(_04376_),
    .X(_04400_));
 sky130_fd_sc_hd__a22o_2 _18489_ (.A1(\alu_shl[7] ),
    .A2(_04400_),
    .B1(_12323_),
    .B2(_04394_),
    .X(_04401_));
 sky130_fd_sc_hd__inv_2 _18490_ (.A(mem_la_wdata[7]),
    .Y(_02336_));
 sky130_fd_sc_hd__o32a_2 _18491_ (.A1(_02336_),
    .A2(_12484_),
    .A3(_04396_),
    .B1(_12322_),
    .B2(_04391_),
    .X(_04402_));
 sky130_vsdinv _18492_ (.A(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__a211o_2 _18493_ (.A1(\alu_shr[7] ),
    .A2(_04399_),
    .B1(_04401_),
    .C1(_04403_),
    .X(_02141_));
 sky130_fd_sc_hd__a22o_2 _18494_ (.A1(\alu_shl[8] ),
    .A2(_04400_),
    .B1(_12348_),
    .B2(_04394_),
    .X(_04404_));
 sky130_fd_sc_hd__inv_2 _18495_ (.A(_11354_),
    .Y(_02339_));
 sky130_fd_sc_hd__o32a_2 _18496_ (.A1(_02339_),
    .A2(_12489_),
    .A3(_04396_),
    .B1(_12347_),
    .B2(_04391_),
    .X(_04405_));
 sky130_vsdinv _18497_ (.A(_04405_),
    .Y(_04406_));
 sky130_fd_sc_hd__a211o_2 _18498_ (.A1(\alu_shr[8] ),
    .A2(_04399_),
    .B1(_04404_),
    .C1(_04406_),
    .X(_02142_));
 sky130_fd_sc_hd__a22o_2 _18499_ (.A1(\alu_shl[9] ),
    .A2(_04400_),
    .B1(_12350_),
    .B2(_04394_),
    .X(_04407_));
 sky130_fd_sc_hd__inv_2 _18500_ (.A(_11353_),
    .Y(_02342_));
 sky130_fd_sc_hd__o32a_2 _18501_ (.A1(_02342_),
    .A2(_12499_),
    .A3(_04396_),
    .B1(_12349_),
    .B2(_04391_),
    .X(_04408_));
 sky130_vsdinv _18502_ (.A(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__a211o_2 _18503_ (.A1(\alu_shr[9] ),
    .A2(_04399_),
    .B1(_04407_),
    .C1(_04409_),
    .X(_02143_));
 sky130_fd_sc_hd__a22o_2 _18504_ (.A1(\alu_shl[10] ),
    .A2(_04400_),
    .B1(_12352_),
    .B2(_04394_),
    .X(_04410_));
 sky130_fd_sc_hd__inv_2 _18505_ (.A(_11352_),
    .Y(_02345_));
 sky130_fd_sc_hd__o32a_2 _18506_ (.A1(_02345_),
    .A2(_12497_),
    .A3(_04396_),
    .B1(_12351_),
    .B2(_04391_),
    .X(_04411_));
 sky130_vsdinv _18507_ (.A(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__a211o_2 _18508_ (.A1(\alu_shr[10] ),
    .A2(_04399_),
    .B1(_04410_),
    .C1(_04412_),
    .X(_02144_));
 sky130_fd_sc_hd__a22o_2 _18509_ (.A1(\alu_shl[11] ),
    .A2(_04400_),
    .B1(_12346_),
    .B2(_04394_),
    .X(_04413_));
 sky130_fd_sc_hd__inv_2 _18510_ (.A(_11351_),
    .Y(_02348_));
 sky130_fd_sc_hd__buf_1 _18511_ (.A(_04364_),
    .X(_04414_));
 sky130_fd_sc_hd__o32a_2 _18512_ (.A1(_02348_),
    .A2(_12503_),
    .A3(_04396_),
    .B1(_12345_),
    .B2(_04414_),
    .X(_04415_));
 sky130_vsdinv _18513_ (.A(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hd__a211o_2 _18514_ (.A1(\alu_shr[11] ),
    .A2(_04399_),
    .B1(_04413_),
    .C1(_04416_),
    .X(_02145_));
 sky130_fd_sc_hd__buf_1 _18515_ (.A(_04358_),
    .X(_04417_));
 sky130_fd_sc_hd__a22o_2 _18516_ (.A1(\alu_shl[12] ),
    .A2(_04400_),
    .B1(_12339_),
    .B2(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__inv_2 _18517_ (.A(_11350_),
    .Y(_02351_));
 sky130_fd_sc_hd__buf_1 _18518_ (.A(_04361_),
    .X(_04419_));
 sky130_fd_sc_hd__o32a_2 _18519_ (.A1(_02351_),
    .A2(_12507_),
    .A3(_04419_),
    .B1(_12338_),
    .B2(_04414_),
    .X(_04420_));
 sky130_vsdinv _18520_ (.A(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__a211o_2 _18521_ (.A1(\alu_shr[12] ),
    .A2(_04399_),
    .B1(_04418_),
    .C1(_04421_),
    .X(_02146_));
 sky130_fd_sc_hd__buf_1 _18522_ (.A(_04369_),
    .X(_04422_));
 sky130_fd_sc_hd__buf_1 _18523_ (.A(_04376_),
    .X(_04423_));
 sky130_fd_sc_hd__a22o_2 _18524_ (.A1(\alu_shl[13] ),
    .A2(_04423_),
    .B1(_12341_),
    .B2(_04417_),
    .X(_04424_));
 sky130_fd_sc_hd__inv_2 _18525_ (.A(_11348_),
    .Y(_02354_));
 sky130_fd_sc_hd__o32a_2 _18526_ (.A1(_02354_),
    .A2(_12512_),
    .A3(_04419_),
    .B1(_12340_),
    .B2(_04414_),
    .X(_04425_));
 sky130_vsdinv _18527_ (.A(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__a211o_2 _18528_ (.A1(\alu_shr[13] ),
    .A2(_04422_),
    .B1(_04424_),
    .C1(_04426_),
    .X(_02147_));
 sky130_fd_sc_hd__a22o_2 _18529_ (.A1(\alu_shl[14] ),
    .A2(_04423_),
    .B1(_12343_),
    .B2(_04417_),
    .X(_04427_));
 sky130_fd_sc_hd__inv_2 _18530_ (.A(_11346_),
    .Y(_02357_));
 sky130_fd_sc_hd__o32a_2 _18531_ (.A1(_02357_),
    .A2(_12516_),
    .A3(_04419_),
    .B1(_12342_),
    .B2(_04414_),
    .X(_04428_));
 sky130_vsdinv _18532_ (.A(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__a211o_2 _18533_ (.A1(\alu_shr[14] ),
    .A2(_04422_),
    .B1(_04427_),
    .C1(_04429_),
    .X(_02148_));
 sky130_fd_sc_hd__a22o_2 _18534_ (.A1(\alu_shl[15] ),
    .A2(_04423_),
    .B1(_12337_),
    .B2(_04417_),
    .X(_04430_));
 sky130_fd_sc_hd__inv_2 _18535_ (.A(_11345_),
    .Y(_02360_));
 sky130_fd_sc_hd__o32a_2 _18536_ (.A1(_02360_),
    .A2(_12520_),
    .A3(_04419_),
    .B1(_12336_),
    .B2(_04414_),
    .X(_04431_));
 sky130_vsdinv _18537_ (.A(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__a211o_2 _18538_ (.A1(\alu_shr[15] ),
    .A2(_04422_),
    .B1(_04430_),
    .C1(_04432_),
    .X(_02149_));
 sky130_fd_sc_hd__a22o_2 _18539_ (.A1(\alu_shl[16] ),
    .A2(_04423_),
    .B1(_12293_),
    .B2(_04417_),
    .X(_04433_));
 sky130_fd_sc_hd__inv_2 _18540_ (.A(pcpi_rs2[16]),
    .Y(_02363_));
 sky130_fd_sc_hd__o32a_2 _18541_ (.A1(_02363_),
    .A2(_12525_),
    .A3(_04419_),
    .B1(_12292_),
    .B2(_04414_),
    .X(_04434_));
 sky130_vsdinv _18542_ (.A(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__a211o_2 _18543_ (.A1(\alu_shr[16] ),
    .A2(_04422_),
    .B1(_04433_),
    .C1(_04435_),
    .X(_02150_));
 sky130_fd_sc_hd__a22o_2 _18544_ (.A1(\alu_shl[17] ),
    .A2(_04423_),
    .B1(_12297_),
    .B2(_04417_),
    .X(_04436_));
 sky130_fd_sc_hd__inv_2 _18545_ (.A(_11344_),
    .Y(_02366_));
 sky130_fd_sc_hd__buf_1 _18546_ (.A(_04363_),
    .X(_04437_));
 sky130_fd_sc_hd__o32a_2 _18547_ (.A1(_02366_),
    .A2(_12536_),
    .A3(_04419_),
    .B1(_12296_),
    .B2(_04437_),
    .X(_04438_));
 sky130_vsdinv _18548_ (.A(_04438_),
    .Y(_04439_));
 sky130_fd_sc_hd__a211o_2 _18549_ (.A1(\alu_shr[17] ),
    .A2(_04422_),
    .B1(_04436_),
    .C1(_04439_),
    .X(_02151_));
 sky130_fd_sc_hd__buf_1 _18550_ (.A(_04358_),
    .X(_04440_));
 sky130_fd_sc_hd__a22o_2 _18551_ (.A1(\alu_shl[18] ),
    .A2(_04423_),
    .B1(_12295_),
    .B2(_04440_),
    .X(_04441_));
 sky130_fd_sc_hd__inv_2 _18552_ (.A(pcpi_rs2[18]),
    .Y(_02369_));
 sky130_fd_sc_hd__buf_1 _18553_ (.A(_04360_),
    .X(_04442_));
 sky130_fd_sc_hd__o32a_2 _18554_ (.A1(_02369_),
    .A2(_12534_),
    .A3(_04442_),
    .B1(_12294_),
    .B2(_04437_),
    .X(_04443_));
 sky130_vsdinv _18555_ (.A(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__a211o_2 _18556_ (.A1(\alu_shr[18] ),
    .A2(_04422_),
    .B1(_04441_),
    .C1(_04444_),
    .X(_02152_));
 sky130_fd_sc_hd__buf_1 _18557_ (.A(_04369_),
    .X(_04445_));
 sky130_fd_sc_hd__buf_1 _18558_ (.A(_04376_),
    .X(_04446_));
 sky130_fd_sc_hd__a22o_2 _18559_ (.A1(\alu_shl[19] ),
    .A2(_04446_),
    .B1(_12299_),
    .B2(_04440_),
    .X(_04447_));
 sky130_fd_sc_hd__inv_2 _18560_ (.A(_11342_),
    .Y(_02372_));
 sky130_fd_sc_hd__o32a_2 _18561_ (.A1(_02372_),
    .A2(_12541_),
    .A3(_04442_),
    .B1(_12298_),
    .B2(_04437_),
    .X(_04448_));
 sky130_vsdinv _18562_ (.A(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__a211o_2 _18563_ (.A1(\alu_shr[19] ),
    .A2(_04445_),
    .B1(_04447_),
    .C1(_04449_),
    .X(_02153_));
 sky130_fd_sc_hd__a22o_2 _18564_ (.A1(\alu_shl[20] ),
    .A2(_04446_),
    .B1(_12290_),
    .B2(_04440_),
    .X(_04450_));
 sky130_fd_sc_hd__inv_2 _18565_ (.A(pcpi_rs2[20]),
    .Y(_02375_));
 sky130_fd_sc_hd__o32a_2 _18566_ (.A1(_02375_),
    .A2(_12545_),
    .A3(_04442_),
    .B1(_12289_),
    .B2(_04437_),
    .X(_04451_));
 sky130_vsdinv _18567_ (.A(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__a211o_2 _18568_ (.A1(\alu_shr[20] ),
    .A2(_04445_),
    .B1(_04450_),
    .C1(_04452_),
    .X(_02154_));
 sky130_fd_sc_hd__a22o_2 _18569_ (.A1(\alu_shl[21] ),
    .A2(_04446_),
    .B1(_12286_),
    .B2(_04440_),
    .X(_04453_));
 sky130_fd_sc_hd__inv_2 _18570_ (.A(_11340_),
    .Y(_02378_));
 sky130_fd_sc_hd__o32a_2 _18571_ (.A1(_02378_),
    .A2(_12549_),
    .A3(_04442_),
    .B1(_12285_),
    .B2(_04437_),
    .X(_04454_));
 sky130_vsdinv _18572_ (.A(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__a211o_2 _18573_ (.A1(\alu_shr[21] ),
    .A2(_04445_),
    .B1(_04453_),
    .C1(_04455_),
    .X(_02155_));
 sky130_fd_sc_hd__a22o_2 _18574_ (.A1(\alu_shl[22] ),
    .A2(_04446_),
    .B1(_12288_),
    .B2(_04440_),
    .X(_04456_));
 sky130_fd_sc_hd__inv_2 _18575_ (.A(pcpi_rs2[22]),
    .Y(_02381_));
 sky130_fd_sc_hd__o32a_2 _18576_ (.A1(_02381_),
    .A2(_12553_),
    .A3(_04442_),
    .B1(_12287_),
    .B2(_04437_),
    .X(_04457_));
 sky130_vsdinv _18577_ (.A(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__a211o_2 _18578_ (.A1(\alu_shr[22] ),
    .A2(_04445_),
    .B1(_04456_),
    .C1(_04458_),
    .X(_02156_));
 sky130_fd_sc_hd__a22o_2 _18579_ (.A1(\alu_shl[23] ),
    .A2(_04446_),
    .B1(_12284_),
    .B2(_04440_),
    .X(_04459_));
 sky130_fd_sc_hd__inv_2 _18580_ (.A(_11339_),
    .Y(_02384_));
 sky130_fd_sc_hd__buf_1 _18581_ (.A(_04363_),
    .X(_04460_));
 sky130_fd_sc_hd__o32a_2 _18582_ (.A1(_02384_),
    .A2(_12557_),
    .A3(_04442_),
    .B1(_12283_),
    .B2(_04460_),
    .X(_04461_));
 sky130_vsdinv _18583_ (.A(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__a211o_2 _18584_ (.A1(\alu_shr[23] ),
    .A2(_04445_),
    .B1(_04459_),
    .C1(_04462_),
    .X(_02157_));
 sky130_fd_sc_hd__buf_1 _18585_ (.A(_04357_),
    .X(_04463_));
 sky130_fd_sc_hd__a22o_2 _18586_ (.A1(\alu_shl[24] ),
    .A2(_04446_),
    .B1(_12317_),
    .B2(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__inv_2 _18587_ (.A(pcpi_rs2[24]),
    .Y(_02387_));
 sky130_fd_sc_hd__buf_1 _18588_ (.A(_04360_),
    .X(_04465_));
 sky130_fd_sc_hd__o32a_2 _18589_ (.A1(_02387_),
    .A2(_12562_),
    .A3(_04465_),
    .B1(_12316_),
    .B2(_04460_),
    .X(_04466_));
 sky130_vsdinv _18590_ (.A(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__a211o_2 _18591_ (.A1(\alu_shr[24] ),
    .A2(_04445_),
    .B1(_04464_),
    .C1(_04467_),
    .X(_02158_));
 sky130_fd_sc_hd__buf_1 _18592_ (.A(_10631_),
    .X(_04468_));
 sky130_fd_sc_hd__buf_1 _18593_ (.A(_04376_),
    .X(_04469_));
 sky130_fd_sc_hd__a22o_2 _18594_ (.A1(\alu_shl[25] ),
    .A2(_04469_),
    .B1(_12315_),
    .B2(_04463_),
    .X(_04470_));
 sky130_fd_sc_hd__inv_2 _18595_ (.A(_11337_),
    .Y(_02390_));
 sky130_fd_sc_hd__o32a_2 _18596_ (.A1(_02390_),
    .A2(_12570_),
    .A3(_04465_),
    .B1(_12314_),
    .B2(_04460_),
    .X(_04471_));
 sky130_vsdinv _18597_ (.A(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hd__a211o_2 _18598_ (.A1(\alu_shr[25] ),
    .A2(_04468_),
    .B1(_04470_),
    .C1(_04472_),
    .X(_02159_));
 sky130_fd_sc_hd__a22o_2 _18599_ (.A1(\alu_shl[26] ),
    .A2(_04469_),
    .B1(_12313_),
    .B2(_04463_),
    .X(_04473_));
 sky130_fd_sc_hd__inv_2 _18600_ (.A(pcpi_rs2[26]),
    .Y(_02393_));
 sky130_fd_sc_hd__o32a_2 _18601_ (.A1(_02393_),
    .A2(_12574_),
    .A3(_04465_),
    .B1(_12312_),
    .B2(_04460_),
    .X(_04474_));
 sky130_vsdinv _18602_ (.A(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__a211o_2 _18603_ (.A1(\alu_shr[26] ),
    .A2(_04468_),
    .B1(_04473_),
    .C1(_04475_),
    .X(_02160_));
 sky130_fd_sc_hd__a22o_2 _18604_ (.A1(\alu_shl[27] ),
    .A2(_04469_),
    .B1(_12311_),
    .B2(_04463_),
    .X(_04476_));
 sky130_fd_sc_hd__inv_2 _18605_ (.A(_11335_),
    .Y(_02396_));
 sky130_fd_sc_hd__o32a_2 _18606_ (.A1(_02396_),
    .A2(_12581_),
    .A3(_04465_),
    .B1(_12310_),
    .B2(_04460_),
    .X(_04477_));
 sky130_vsdinv _18607_ (.A(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__a211o_2 _18608_ (.A1(\alu_shr[27] ),
    .A2(_04468_),
    .B1(_04476_),
    .C1(_04478_),
    .X(_02161_));
 sky130_fd_sc_hd__a22o_2 _18609_ (.A1(\alu_shl[28] ),
    .A2(_04469_),
    .B1(_12304_),
    .B2(_04463_),
    .X(_04479_));
 sky130_fd_sc_hd__inv_2 _18610_ (.A(pcpi_rs2[28]),
    .Y(_02399_));
 sky130_fd_sc_hd__o32a_2 _18611_ (.A1(_02399_),
    .A2(_12590_),
    .A3(_04465_),
    .B1(_12303_),
    .B2(_04460_),
    .X(_04480_));
 sky130_vsdinv _18612_ (.A(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__a211o_2 _18613_ (.A1(\alu_shr[28] ),
    .A2(_04468_),
    .B1(_04479_),
    .C1(_04481_),
    .X(_02162_));
 sky130_fd_sc_hd__a22o_2 _18614_ (.A1(\alu_shl[29] ),
    .A2(_04469_),
    .B1(_12302_),
    .B2(_04463_),
    .X(_04482_));
 sky130_fd_sc_hd__inv_2 _18615_ (.A(_11334_),
    .Y(_02402_));
 sky130_fd_sc_hd__o32a_2 _18616_ (.A1(_02402_),
    .A2(_12597_),
    .A3(_04465_),
    .B1(_12301_),
    .B2(_04364_),
    .X(_04483_));
 sky130_vsdinv _18617_ (.A(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__a211o_2 _18618_ (.A1(\alu_shr[29] ),
    .A2(_04468_),
    .B1(_04482_),
    .C1(_04484_),
    .X(_02163_));
 sky130_fd_sc_hd__a22o_2 _18619_ (.A1(\alu_shl[30] ),
    .A2(_04469_),
    .B1(_12308_),
    .B2(_04358_),
    .X(_04485_));
 sky130_fd_sc_hd__inv_2 _18620_ (.A(pcpi_rs2[30]),
    .Y(_02405_));
 sky130_fd_sc_hd__o32a_2 _18621_ (.A1(_02405_),
    .A2(_12595_),
    .A3(_04361_),
    .B1(_12307_),
    .B2(_04364_),
    .X(_04486_));
 sky130_vsdinv _18622_ (.A(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__a211o_2 _18623_ (.A1(\alu_shr[30] ),
    .A2(_04468_),
    .B1(_04485_),
    .C1(_04487_),
    .X(_02164_));
 sky130_fd_sc_hd__a22o_2 _18624_ (.A1(\alu_shl[31] ),
    .A2(_04376_),
    .B1(_12306_),
    .B2(_04358_),
    .X(_04488_));
 sky130_fd_sc_hd__o32a_2 _18625_ (.A1(_10568_),
    .A2(_10594_),
    .A3(_04361_),
    .B1(_12305_),
    .B2(_04364_),
    .X(_04489_));
 sky130_vsdinv _18626_ (.A(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__a211o_2 _18627_ (.A1(\alu_shr[31] ),
    .A2(_04369_),
    .B1(_04488_),
    .C1(_04490_),
    .X(_02165_));
 sky130_fd_sc_hd__and3_2 _18628_ (.A(_10490_),
    .B(_10811_),
    .C(_00289_),
    .X(_02166_));
 sky130_vsdinv _18629_ (.A(_12773_),
    .Y(mem_la_wstrb[1]));
 sky130_vsdinv _18630_ (.A(_12776_),
    .Y(mem_la_wstrb[2]));
 sky130_vsdinv _18631_ (.A(_12778_),
    .Y(mem_la_wstrb[3]));
 sky130_fd_sc_hd__buf_1 _18632_ (.A(\mem_wordsize[1] ),
    .X(_04491_));
 sky130_fd_sc_hd__a22o_2 _18633_ (.A1(_11364_),
    .A2(_04491_),
    .B1(_11354_),
    .B2(_04100_),
    .X(_02167_));
 sky130_fd_sc_hd__a22o_2 _18634_ (.A1(_11363_),
    .A2(_04491_),
    .B1(_11353_),
    .B2(_04100_),
    .X(_02168_));
 sky130_fd_sc_hd__a22o_2 _18635_ (.A1(_11362_),
    .A2(_04491_),
    .B1(_11352_),
    .B2(_04100_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_2 _18636_ (.A1(_11361_),
    .A2(_04491_),
    .B1(_11351_),
    .B2(_04100_),
    .X(_02170_));
 sky130_fd_sc_hd__a22o_2 _18637_ (.A1(_11360_),
    .A2(_04491_),
    .B1(_11350_),
    .B2(_12901_),
    .X(_02171_));
 sky130_fd_sc_hd__a22o_2 _18638_ (.A1(_11359_),
    .A2(_04491_),
    .B1(_11348_),
    .B2(_12901_),
    .X(_02172_));
 sky130_fd_sc_hd__a22o_2 _18639_ (.A1(_11358_),
    .A2(\mem_wordsize[1] ),
    .B1(_11346_),
    .B2(_12901_),
    .X(_02173_));
 sky130_fd_sc_hd__a22o_2 _18640_ (.A1(_11356_),
    .A2(\mem_wordsize[1] ),
    .B1(_11345_),
    .B2(_12901_),
    .X(_02174_));
 sky130_fd_sc_hd__nor2_2 _18641_ (.A(_12281_),
    .B(_01683_),
    .Y(_02175_));
 sky130_fd_sc_hd__nor2_2 _18642_ (.A(_02318_),
    .B(_01683_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_2 _18643_ (.A(_02321_),
    .B(_01683_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_2 _18644_ (.A(_02324_),
    .B(_01683_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_2 _18645_ (.A(_02327_),
    .B(_01683_),
    .Y(_02179_));
 sky130_fd_sc_hd__nor2_2 _18646_ (.A(_02330_),
    .B(_12769_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_2 _18647_ (.A(_02333_),
    .B(_12769_),
    .Y(_02181_));
 sky130_fd_sc_hd__nor2_2 _18648_ (.A(_02336_),
    .B(_12769_),
    .Y(_02182_));
 sky130_fd_sc_hd__or2_2 _18649_ (.A(_11255_),
    .B(_11256_),
    .X(_02183_));
 sky130_fd_sc_hd__or2_2 _18650_ (.A(\irq_pending[3] ),
    .B(irq[3]),
    .X(_02214_));
 sky130_fd_sc_hd__and2_2 _18651_ (.A(\irq_mask[3] ),
    .B(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__or2_2 _18652_ (.A(\irq_pending[4] ),
    .B(irq[4]),
    .X(_02218_));
 sky130_fd_sc_hd__and2_2 _18653_ (.A(\irq_mask[4] ),
    .B(_02218_),
    .X(_02219_));
 sky130_fd_sc_hd__or2_2 _18654_ (.A(\irq_pending[5] ),
    .B(irq[5]),
    .X(_02221_));
 sky130_fd_sc_hd__and2_2 _18655_ (.A(\irq_mask[5] ),
    .B(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__or2_2 _18656_ (.A(\irq_pending[6] ),
    .B(irq[6]),
    .X(_02224_));
 sky130_fd_sc_hd__and2_2 _18657_ (.A(\irq_mask[6] ),
    .B(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__or2_2 _18658_ (.A(\irq_pending[7] ),
    .B(irq[7]),
    .X(_02227_));
 sky130_fd_sc_hd__and2_2 _18659_ (.A(\irq_mask[7] ),
    .B(_02227_),
    .X(_02228_));
 sky130_fd_sc_hd__or2_2 _18660_ (.A(\irq_pending[8] ),
    .B(irq[8]),
    .X(_02230_));
 sky130_fd_sc_hd__and2_2 _18661_ (.A(\irq_mask[8] ),
    .B(_02230_),
    .X(_02231_));
 sky130_fd_sc_hd__or2_2 _18662_ (.A(\irq_pending[9] ),
    .B(irq[9]),
    .X(_02233_));
 sky130_fd_sc_hd__and2_2 _18663_ (.A(\irq_mask[9] ),
    .B(_02233_),
    .X(_02234_));
 sky130_fd_sc_hd__or2_2 _18664_ (.A(\irq_pending[10] ),
    .B(irq[10]),
    .X(_02236_));
 sky130_fd_sc_hd__and2_2 _18665_ (.A(\irq_mask[10] ),
    .B(_02236_),
    .X(_02237_));
 sky130_fd_sc_hd__or2_2 _18666_ (.A(\irq_pending[11] ),
    .B(irq[11]),
    .X(_02239_));
 sky130_fd_sc_hd__and2_2 _18667_ (.A(\irq_mask[11] ),
    .B(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__or2_2 _18668_ (.A(\irq_pending[12] ),
    .B(irq[12]),
    .X(_02242_));
 sky130_fd_sc_hd__and2_2 _18669_ (.A(\irq_mask[12] ),
    .B(_02242_),
    .X(_02243_));
 sky130_fd_sc_hd__or2_2 _18670_ (.A(\irq_pending[13] ),
    .B(irq[13]),
    .X(_02245_));
 sky130_fd_sc_hd__and2_2 _18671_ (.A(\irq_mask[13] ),
    .B(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__or2_2 _18672_ (.A(\irq_pending[14] ),
    .B(irq[14]),
    .X(_02248_));
 sky130_fd_sc_hd__and2_2 _18673_ (.A(\irq_mask[14] ),
    .B(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__or2_2 _18674_ (.A(\irq_pending[15] ),
    .B(irq[15]),
    .X(_02251_));
 sky130_fd_sc_hd__and2_2 _18675_ (.A(\irq_mask[15] ),
    .B(_02251_),
    .X(_02252_));
 sky130_fd_sc_hd__or2_2 _18676_ (.A(\irq_pending[16] ),
    .B(irq[16]),
    .X(_02254_));
 sky130_fd_sc_hd__and2_2 _18677_ (.A(\irq_mask[16] ),
    .B(_02254_),
    .X(_02255_));
 sky130_fd_sc_hd__or2_2 _18678_ (.A(\irq_pending[17] ),
    .B(irq[17]),
    .X(_02257_));
 sky130_fd_sc_hd__and2_2 _18679_ (.A(\irq_mask[17] ),
    .B(_02257_),
    .X(_02258_));
 sky130_fd_sc_hd__or2_2 _18680_ (.A(\irq_pending[18] ),
    .B(irq[18]),
    .X(_02260_));
 sky130_fd_sc_hd__and2_2 _18681_ (.A(\irq_mask[18] ),
    .B(_02260_),
    .X(_02261_));
 sky130_fd_sc_hd__or2_2 _18682_ (.A(\irq_pending[19] ),
    .B(irq[19]),
    .X(_02263_));
 sky130_fd_sc_hd__and2_2 _18683_ (.A(\irq_mask[19] ),
    .B(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__or2_2 _18684_ (.A(\irq_pending[20] ),
    .B(irq[20]),
    .X(_02266_));
 sky130_fd_sc_hd__and2_2 _18685_ (.A(\irq_mask[20] ),
    .B(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__or2_2 _18686_ (.A(\irq_pending[21] ),
    .B(irq[21]),
    .X(_02269_));
 sky130_fd_sc_hd__and2_2 _18687_ (.A(\irq_mask[21] ),
    .B(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__or2_2 _18688_ (.A(\irq_pending[22] ),
    .B(irq[22]),
    .X(_02272_));
 sky130_fd_sc_hd__and2_2 _18689_ (.A(\irq_mask[22] ),
    .B(_02272_),
    .X(_02273_));
 sky130_fd_sc_hd__or2_2 _18690_ (.A(\irq_pending[23] ),
    .B(irq[23]),
    .X(_02275_));
 sky130_fd_sc_hd__and2_2 _18691_ (.A(\irq_mask[23] ),
    .B(_02275_),
    .X(_02276_));
 sky130_fd_sc_hd__or2_2 _18692_ (.A(\irq_pending[24] ),
    .B(irq[24]),
    .X(_02278_));
 sky130_fd_sc_hd__and2_2 _18693_ (.A(\irq_mask[24] ),
    .B(_02278_),
    .X(_02279_));
 sky130_fd_sc_hd__or2_2 _18694_ (.A(\irq_pending[25] ),
    .B(irq[25]),
    .X(_02281_));
 sky130_fd_sc_hd__and2_2 _18695_ (.A(\irq_mask[25] ),
    .B(_02281_),
    .X(_02282_));
 sky130_fd_sc_hd__or2_2 _18696_ (.A(\irq_pending[26] ),
    .B(irq[26]),
    .X(_02284_));
 sky130_fd_sc_hd__and2_2 _18697_ (.A(\irq_mask[26] ),
    .B(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__or2_2 _18698_ (.A(\irq_pending[27] ),
    .B(irq[27]),
    .X(_02287_));
 sky130_fd_sc_hd__and2_2 _18699_ (.A(\irq_mask[27] ),
    .B(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__or2_2 _18700_ (.A(\irq_pending[28] ),
    .B(irq[28]),
    .X(_02290_));
 sky130_fd_sc_hd__and2_2 _18701_ (.A(\irq_mask[28] ),
    .B(_02290_),
    .X(_02291_));
 sky130_fd_sc_hd__or2_2 _18702_ (.A(\irq_pending[29] ),
    .B(irq[29]),
    .X(_02293_));
 sky130_fd_sc_hd__and2_2 _18703_ (.A(\irq_mask[29] ),
    .B(_02293_),
    .X(_02294_));
 sky130_fd_sc_hd__or2_2 _18704_ (.A(\irq_pending[30] ),
    .B(irq[30]),
    .X(_02296_));
 sky130_fd_sc_hd__and2_2 _18705_ (.A(\irq_mask[30] ),
    .B(_02296_),
    .X(_02297_));
 sky130_fd_sc_hd__or2_2 _18706_ (.A(\irq_pending[31] ),
    .B(irq[31]),
    .X(_02299_));
 sky130_fd_sc_hd__and2_2 _18707_ (.A(\irq_mask[31] ),
    .B(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__or4_2 _18708_ (.A(\timer[3] ),
    .B(\timer[2] ),
    .C(\timer[7] ),
    .D(\timer[6] ),
    .X(_04492_));
 sky130_fd_sc_hd__or4_2 _18709_ (.A(\timer[19] ),
    .B(\timer[18] ),
    .C(\timer[15] ),
    .D(\timer[14] ),
    .X(_04493_));
 sky130_fd_sc_hd__or4_2 _18710_ (.A(\timer[21] ),
    .B(\timer[20] ),
    .C(\timer[23] ),
    .D(\timer[22] ),
    .X(_04494_));
 sky130_fd_sc_hd__or4_2 _18711_ (.A(\timer[31] ),
    .B(\timer[30] ),
    .C(\timer[27] ),
    .D(\timer[26] ),
    .X(_04495_));
 sky130_fd_sc_hd__or4_2 _18712_ (.A(_04492_),
    .B(_04493_),
    .C(_04494_),
    .D(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__or4_2 _18713_ (.A(\timer[9] ),
    .B(\timer[8] ),
    .C(\timer[11] ),
    .D(\timer[10] ),
    .X(_04497_));
 sky130_fd_sc_hd__or4_2 _18714_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .C(\timer[29] ),
    .D(\timer[28] ),
    .X(_04498_));
 sky130_fd_sc_hd__or4_2 _18715_ (.A(\timer[25] ),
    .B(\timer[24] ),
    .C(\timer[1] ),
    .D(_12409_),
    .X(_04499_));
 sky130_fd_sc_hd__or4_2 _18716_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .C(\timer[17] ),
    .D(\timer[16] ),
    .X(_04500_));
 sky130_fd_sc_hd__or4_2 _18717_ (.A(_04497_),
    .B(_04498_),
    .C(_04499_),
    .D(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__o21ai_2 _18718_ (.A1(_04496_),
    .A2(_04501_),
    .B1(_10512_),
    .Y(_02302_));
 sky130_fd_sc_hd__or2_2 _18719_ (.A(_02303_),
    .B(irq[0]),
    .X(_02304_));
 sky130_fd_sc_hd__and2_2 _18720_ (.A(\irq_mask[0] ),
    .B(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__nor2_2 _18721_ (.A(\irq_pending[2] ),
    .B(irq[2]),
    .Y(_02307_));
 sky130_fd_sc_hd__or2_2 _18722_ (.A(_10511_),
    .B(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__nor2_2 _18723_ (.A(_10688_),
    .B(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__or2_2 _18724_ (.A(_12226_),
    .B(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__or2_2 _18725_ (.A(_02313_),
    .B(_12226_),
    .X(_02314_));
 sky130_fd_sc_hd__or2_2 _18726_ (.A(_02316_),
    .B(_12226_),
    .X(_02317_));
 sky130_fd_sc_hd__o32a_2 _18727_ (.A1(_02387_),
    .A2(pcpi_rs1[24]),
    .A3(_12315_),
    .B1(_02390_),
    .B2(_11824_),
    .X(_04502_));
 sky130_fd_sc_hd__o22a_2 _18728_ (.A1(_02393_),
    .A2(_11821_),
    .B1(_12313_),
    .B2(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__o22a_2 _18729_ (.A1(_02396_),
    .A2(_11819_),
    .B1(_12311_),
    .B2(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__o22a_2 _18730_ (.A1(_02399_),
    .A2(pcpi_rs1[28]),
    .B1(_12304_),
    .B2(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__o22a_2 _18731_ (.A1(_02402_),
    .A2(pcpi_rs1[29]),
    .B1(_12302_),
    .B2(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__or2_2 _18732_ (.A(_12309_),
    .B(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__o32a_2 _18733_ (.A1(_02363_),
    .A2(_11839_),
    .A3(_12297_),
    .B1(_02366_),
    .B2(_11838_),
    .X(_04508_));
 sky130_fd_sc_hd__o22a_2 _18734_ (.A1(_02369_),
    .A2(_11836_),
    .B1(_12295_),
    .B2(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__o22a_2 _18735_ (.A1(_02372_),
    .A2(_11834_),
    .B1(_12299_),
    .B2(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__o22a_2 _18736_ (.A1(_02375_),
    .A2(_11832_),
    .B1(_12290_),
    .B2(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__o22a_2 _18737_ (.A1(_02378_),
    .A2(_11831_),
    .B1(_12286_),
    .B2(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__o22a_2 _18738_ (.A1(_02381_),
    .A2(_11830_),
    .B1(_12288_),
    .B2(_04512_),
    .X(_04513_));
 sky130_fd_sc_hd__o32a_2 _18739_ (.A1(_02351_),
    .A2(_11845_),
    .A3(_12341_),
    .B1(_02354_),
    .B2(_11843_),
    .X(_04514_));
 sky130_fd_sc_hd__o22a_2 _18740_ (.A1(_02357_),
    .A2(_11841_),
    .B1(_12343_),
    .B2(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__o21a_2 _18741_ (.A1(_12192_),
    .A2(_00048_),
    .B1(_11861_),
    .X(_04516_));
 sky130_fd_sc_hd__o32a_2 _18742_ (.A1(_00049_),
    .A2(_12334_),
    .A3(_04516_),
    .B1(_12191_),
    .B2(_11860_),
    .X(_04517_));
 sky130_fd_sc_hd__o22a_2 _18743_ (.A1(_12187_),
    .A2(_11859_),
    .B1(_12327_),
    .B2(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__o22a_2 _18744_ (.A1(_12185_),
    .A2(_11858_),
    .B1(_12330_),
    .B2(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__o22a_2 _18745_ (.A1(_02330_),
    .A2(_11857_),
    .B1(_12321_),
    .B2(_04519_),
    .X(_04520_));
 sky130_fd_sc_hd__o22a_2 _18746_ (.A1(_02333_),
    .A2(_11856_),
    .B1(_12332_),
    .B2(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__o22a_2 _18747_ (.A1(_02336_),
    .A2(_11853_),
    .B1(_12323_),
    .B2(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__o32a_2 _18748_ (.A1(_02339_),
    .A2(_11850_),
    .A3(_12350_),
    .B1(_02342_),
    .B2(_11849_),
    .X(_04523_));
 sky130_fd_sc_hd__o22a_2 _18749_ (.A1(_02345_),
    .A2(_11847_),
    .B1(_12352_),
    .B2(_04523_),
    .X(_04524_));
 sky130_fd_sc_hd__or2_2 _18750_ (.A(_12346_),
    .B(_04524_),
    .X(_04525_));
 sky130_fd_sc_hd__o221a_2 _18751_ (.A1(_02348_),
    .A2(_11846_),
    .B1(_12353_),
    .B2(_04522_),
    .C1(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__or2_2 _18752_ (.A(_12344_),
    .B(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__o221ai_2 _18753_ (.A1(_02360_),
    .A2(_11840_),
    .B1(_12337_),
    .B2(_04515_),
    .C1(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__or3b_2 _18754_ (.A(_12291_),
    .B(_12300_),
    .C_N(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__o221a_2 _18755_ (.A1(_02384_),
    .A2(_11829_),
    .B1(_12284_),
    .B2(_04513_),
    .C1(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__or2_2 _18756_ (.A(_12319_),
    .B(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__o311a_2 _18757_ (.A1(_02405_),
    .A2(_11816_),
    .A3(_12306_),
    .B1(_04507_),
    .C1(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__o21a_2 _18758_ (.A1(_11812_),
    .A2(_10594_),
    .B1(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__nor2_2 _18759_ (.A(_00000_),
    .B(_04533_),
    .Y(_00002_));
 sky130_vsdinv _18760_ (.A(_04532_),
    .Y(_04534_));
 sky130_fd_sc_hd__o221a_2 _18761_ (.A1(_12306_),
    .A2(_04534_),
    .B1(_11812_),
    .B2(_10594_),
    .C1(_12355_),
    .X(_00001_));
 sky130_vsdinv _18762_ (.A(\pcpi_mul.rs2[0] ),
    .Y(_04535_));
 sky130_fd_sc_hd__buf_1 _18763_ (.A(_04535_),
    .X(_04536_));
 sky130_fd_sc_hd__buf_1 _18764_ (.A(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__buf_1 _18765_ (.A(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__buf_1 _18766_ (.A(_04538_),
    .X(_04539_));
 sky130_vsdinv _18767_ (.A(\pcpi_mul.rs1[0] ),
    .Y(_04540_));
 sky130_fd_sc_hd__buf_1 _18768_ (.A(_04540_),
    .X(_04541_));
 sky130_fd_sc_hd__buf_1 _18769_ (.A(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__buf_1 _18770_ (.A(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__buf_1 _18771_ (.A(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__buf_1 _18772_ (.A(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__buf_1 _18773_ (.A(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__nor2_2 _18774_ (.A(_04539_),
    .B(_04546_),
    .Y(_02623_));
 sky130_fd_sc_hd__or2_2 _18775_ (.A(mem_la_wdata[1]),
    .B(mem_la_wdata[0]),
    .X(_04547_));
 sky130_fd_sc_hd__o21ai_2 _18776_ (.A1(_02318_),
    .A2(_12281_),
    .B1(_04547_),
    .Y(_02319_));
 sky130_vsdinv _18777_ (.A(_02320_),
    .Y(_04548_));
 sky130_fd_sc_hd__o22a_2 _18778_ (.A1(_12451_),
    .A2(_04548_),
    .B1(_11861_),
    .B2(_02320_),
    .X(_04549_));
 sky130_vsdinv _18779_ (.A(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__o32a_2 _18780_ (.A1(_12281_),
    .A2(_11863_),
    .A3(_04549_),
    .B1(_12282_),
    .B2(_04550_),
    .X(_02602_));
 sky130_fd_sc_hd__or2_2 _18781_ (.A(mem_la_wdata[2]),
    .B(_04547_),
    .X(_04551_));
 sky130_fd_sc_hd__a21bo_2 _18782_ (.A1(_11362_),
    .A2(_04547_),
    .B1_N(_04551_),
    .X(_02322_));
 sky130_fd_sc_hd__o22a_2 _18783_ (.A1(_12451_),
    .A2(_04548_),
    .B1(_12282_),
    .B2(_04550_),
    .X(_04552_));
 sky130_fd_sc_hd__nor2_2 _18784_ (.A(pcpi_rs1[2]),
    .B(_02323_),
    .Y(_04553_));
 sky130_fd_sc_hd__a21o_2 _18785_ (.A1(_11860_),
    .A2(_02323_),
    .B1(_04553_),
    .X(_04554_));
 sky130_fd_sc_hd__o2bb2a_2 _18786_ (.A1_N(_04552_),
    .A2_N(_04554_),
    .B1(_04552_),
    .B2(_04554_),
    .X(_02613_));
 sky130_fd_sc_hd__or2_2 _18787_ (.A(mem_la_wdata[3]),
    .B(_04551_),
    .X(_04555_));
 sky130_vsdinv _18788_ (.A(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__a21o_2 _18789_ (.A1(_11361_),
    .A2(_04551_),
    .B1(_04556_),
    .X(_02325_));
 sky130_fd_sc_hd__o2bb2a_2 _18790_ (.A1_N(pcpi_rs1[2]),
    .A2_N(_02323_),
    .B1(_04552_),
    .B2(_04553_),
    .X(_04557_));
 sky130_fd_sc_hd__nor2_2 _18791_ (.A(pcpi_rs1[3]),
    .B(_02326_),
    .Y(_04558_));
 sky130_fd_sc_hd__a21o_2 _18792_ (.A1(_11859_),
    .A2(_02326_),
    .B1(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__o2bb2a_2 _18793_ (.A1_N(_04557_),
    .A2_N(_04559_),
    .B1(_04557_),
    .B2(_04559_),
    .X(_02616_));
 sky130_fd_sc_hd__or2_2 _18794_ (.A(mem_la_wdata[4]),
    .B(_04555_),
    .X(_04560_));
 sky130_fd_sc_hd__o21ai_2 _18795_ (.A1(_02327_),
    .A2(_04556_),
    .B1(_04560_),
    .Y(_02328_));
 sky130_fd_sc_hd__o2bb2a_2 _18796_ (.A1_N(pcpi_rs1[3]),
    .A2_N(_02326_),
    .B1(_04557_),
    .B2(_04558_),
    .X(_04561_));
 sky130_fd_sc_hd__nor2_2 _18797_ (.A(pcpi_rs1[4]),
    .B(_02329_),
    .Y(_04562_));
 sky130_fd_sc_hd__a21o_2 _18798_ (.A1(_11858_),
    .A2(_02329_),
    .B1(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__o2bb2a_2 _18799_ (.A1_N(_04561_),
    .A2_N(_04563_),
    .B1(_04561_),
    .B2(_04563_),
    .X(_02617_));
 sky130_fd_sc_hd__or2_2 _18800_ (.A(mem_la_wdata[5]),
    .B(_04560_),
    .X(_04564_));
 sky130_vsdinv _18801_ (.A(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__a21o_2 _18802_ (.A1(_11359_),
    .A2(_04560_),
    .B1(_04565_),
    .X(_02331_));
 sky130_fd_sc_hd__o2bb2a_2 _18803_ (.A1_N(pcpi_rs1[4]),
    .A2_N(_02329_),
    .B1(_04561_),
    .B2(_04562_),
    .X(_04566_));
 sky130_fd_sc_hd__nor2_2 _18804_ (.A(pcpi_rs1[5]),
    .B(_02332_),
    .Y(_04567_));
 sky130_fd_sc_hd__a21o_2 _18805_ (.A1(_11857_),
    .A2(_02332_),
    .B1(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__o2bb2a_2 _18806_ (.A1_N(_04566_),
    .A2_N(_04568_),
    .B1(_04566_),
    .B2(_04568_),
    .X(_02618_));
 sky130_fd_sc_hd__or2_2 _18807_ (.A(mem_la_wdata[6]),
    .B(_04564_),
    .X(_04569_));
 sky130_fd_sc_hd__o21ai_2 _18808_ (.A1(_02333_),
    .A2(_04565_),
    .B1(_04569_),
    .Y(_02334_));
 sky130_fd_sc_hd__o2bb2ai_2 _18809_ (.A1_N(pcpi_rs1[5]),
    .A2_N(_02332_),
    .B1(_04566_),
    .B2(_04567_),
    .Y(_04570_));
 sky130_fd_sc_hd__o2bb2a_2 _18810_ (.A1_N(_11855_),
    .A2_N(_02335_),
    .B1(_11855_),
    .B2(_02335_),
    .X(_04571_));
 sky130_fd_sc_hd__o2bb2a_2 _18811_ (.A1_N(_04570_),
    .A2_N(_04571_),
    .B1(_04570_),
    .B2(_04571_),
    .X(_02619_));
 sky130_fd_sc_hd__or2_2 _18812_ (.A(mem_la_wdata[7]),
    .B(_04569_),
    .X(_04572_));
 sky130_vsdinv _18813_ (.A(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__a21o_2 _18814_ (.A1(_11356_),
    .A2(_04569_),
    .B1(_04573_),
    .X(_02337_));
 sky130_fd_sc_hd__o2bb2a_2 _18815_ (.A1_N(_11852_),
    .A2_N(_02338_),
    .B1(_11852_),
    .B2(_02338_),
    .X(_04574_));
 sky130_fd_sc_hd__a22o_2 _18816_ (.A1(_11856_),
    .A2(_02335_),
    .B1(_04570_),
    .B2(_04571_),
    .X(_04575_));
 sky130_fd_sc_hd__a2bb2oi_2 _18817_ (.A1_N(_04574_),
    .A2_N(_04575_),
    .B1(_04574_),
    .B2(_04575_),
    .Y(_02620_));
 sky130_fd_sc_hd__or2_2 _18818_ (.A(pcpi_rs2[8]),
    .B(_04572_),
    .X(_04576_));
 sky130_fd_sc_hd__o21ai_2 _18819_ (.A1(_02339_),
    .A2(_04573_),
    .B1(_04576_),
    .Y(_02340_));
 sky130_fd_sc_hd__or2_2 _18820_ (.A(_11852_),
    .B(_02338_),
    .X(_04577_));
 sky130_fd_sc_hd__a32o_2 _18821_ (.A1(_11855_),
    .A2(_02335_),
    .A3(_04577_),
    .B1(_11853_),
    .B2(_02338_),
    .X(_04578_));
 sky130_fd_sc_hd__a31o_2 _18822_ (.A1(_04571_),
    .A2(_04574_),
    .A3(_04570_),
    .B1(_04578_),
    .X(_04579_));
 sky130_fd_sc_hd__o2bb2a_2 _18823_ (.A1_N(pcpi_rs1[8]),
    .A2_N(_02341_),
    .B1(pcpi_rs1[8]),
    .B2(_02341_),
    .X(_04580_));
 sky130_fd_sc_hd__o2bb2a_2 _18824_ (.A1_N(_04579_),
    .A2_N(_04580_),
    .B1(_04579_),
    .B2(_04580_),
    .X(_02621_));
 sky130_fd_sc_hd__or2_2 _18825_ (.A(pcpi_rs2[9]),
    .B(_04576_),
    .X(_04581_));
 sky130_vsdinv _18826_ (.A(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__a21o_2 _18827_ (.A1(_11353_),
    .A2(_04576_),
    .B1(_04582_),
    .X(_02343_));
 sky130_fd_sc_hd__o2bb2a_2 _18828_ (.A1_N(_11848_),
    .A2_N(_02344_),
    .B1(_11848_),
    .B2(_02344_),
    .X(_04583_));
 sky130_fd_sc_hd__a22o_2 _18829_ (.A1(_11850_),
    .A2(_02341_),
    .B1(_04579_),
    .B2(_04580_),
    .X(_04584_));
 sky130_fd_sc_hd__a2bb2oi_2 _18830_ (.A1_N(_04583_),
    .A2_N(_04584_),
    .B1(_04583_),
    .B2(_04584_),
    .Y(_02622_));
 sky130_fd_sc_hd__or2_2 _18831_ (.A(pcpi_rs2[10]),
    .B(_04581_),
    .X(_04585_));
 sky130_fd_sc_hd__o21ai_2 _18832_ (.A1(_02345_),
    .A2(_04582_),
    .B1(_04585_),
    .Y(_02346_));
 sky130_vsdinv _18833_ (.A(_02347_),
    .Y(_04586_));
 sky130_fd_sc_hd__a22o_2 _18834_ (.A1(_11847_),
    .A2(_02347_),
    .B1(_12497_),
    .B2(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__or2_2 _18835_ (.A(pcpi_rs1[9]),
    .B(_02344_),
    .X(_04588_));
 sky130_fd_sc_hd__a32o_2 _18836_ (.A1(pcpi_rs1[8]),
    .A2(_02341_),
    .A3(_04588_),
    .B1(_11849_),
    .B2(_02344_),
    .X(_04589_));
 sky130_fd_sc_hd__a31oi_2 _18837_ (.A1(_04580_),
    .A2(_04583_),
    .A3(_04579_),
    .B1(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__a2bb2oi_2 _18838_ (.A1_N(_04587_),
    .A2_N(_04590_),
    .B1(_04587_),
    .B2(_04590_),
    .Y(_02592_));
 sky130_fd_sc_hd__or2_2 _18839_ (.A(pcpi_rs2[11]),
    .B(_04585_),
    .X(_04591_));
 sky130_vsdinv _18840_ (.A(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__a21o_2 _18841_ (.A1(_11351_),
    .A2(_04585_),
    .B1(_04592_),
    .X(_02349_));
 sky130_vsdinv _18842_ (.A(_02350_),
    .Y(_04593_));
 sky130_fd_sc_hd__a22o_2 _18843_ (.A1(_11846_),
    .A2(_02350_),
    .B1(_12503_),
    .B2(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__o22a_2 _18844_ (.A1(_12497_),
    .A2(_04586_),
    .B1(_04587_),
    .B2(_04590_),
    .X(_04595_));
 sky130_fd_sc_hd__a2bb2oi_2 _18845_ (.A1_N(_04594_),
    .A2_N(_04595_),
    .B1(_04594_),
    .B2(_04595_),
    .Y(_02593_));
 sky130_fd_sc_hd__or2_2 _18846_ (.A(pcpi_rs2[12]),
    .B(_04591_),
    .X(_04596_));
 sky130_fd_sc_hd__o21ai_2 _18847_ (.A1(_02351_),
    .A2(_04592_),
    .B1(_04596_),
    .Y(_02352_));
 sky130_vsdinv _18848_ (.A(_02353_),
    .Y(_04597_));
 sky130_fd_sc_hd__a22o_2 _18849_ (.A1(_11845_),
    .A2(_02353_),
    .B1(_12507_),
    .B2(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__o22a_2 _18850_ (.A1(_12503_),
    .A2(_04593_),
    .B1(_04594_),
    .B2(_04595_),
    .X(_04599_));
 sky130_fd_sc_hd__a2bb2oi_2 _18851_ (.A1_N(_04598_),
    .A2_N(_04599_),
    .B1(_04598_),
    .B2(_04599_),
    .Y(_02594_));
 sky130_fd_sc_hd__or2_2 _18852_ (.A(pcpi_rs2[13]),
    .B(_04596_),
    .X(_04600_));
 sky130_vsdinv _18853_ (.A(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__a21o_2 _18854_ (.A1(_11348_),
    .A2(_04596_),
    .B1(_04601_),
    .X(_02355_));
 sky130_vsdinv _18855_ (.A(_02356_),
    .Y(_04602_));
 sky130_fd_sc_hd__a22o_2 _18856_ (.A1(_11843_),
    .A2(_02356_),
    .B1(_12512_),
    .B2(_04602_),
    .X(_04603_));
 sky130_fd_sc_hd__o22a_2 _18857_ (.A1(_12507_),
    .A2(_04597_),
    .B1(_04598_),
    .B2(_04599_),
    .X(_04604_));
 sky130_fd_sc_hd__a2bb2oi_2 _18858_ (.A1_N(_04603_),
    .A2_N(_04604_),
    .B1(_04603_),
    .B2(_04604_),
    .Y(_02595_));
 sky130_fd_sc_hd__or2_2 _18859_ (.A(pcpi_rs2[14]),
    .B(_04600_),
    .X(_04605_));
 sky130_fd_sc_hd__o21ai_2 _18860_ (.A1(_02357_),
    .A2(_04601_),
    .B1(_04605_),
    .Y(_02358_));
 sky130_vsdinv _18861_ (.A(_02359_),
    .Y(_04606_));
 sky130_fd_sc_hd__a22o_2 _18862_ (.A1(_11841_),
    .A2(_02359_),
    .B1(_12516_),
    .B2(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__o22a_2 _18863_ (.A1(_12512_),
    .A2(_04602_),
    .B1(_04603_),
    .B2(_04604_),
    .X(_04608_));
 sky130_fd_sc_hd__a2bb2oi_2 _18864_ (.A1_N(_04607_),
    .A2_N(_04608_),
    .B1(_04607_),
    .B2(_04608_),
    .Y(_02596_));
 sky130_fd_sc_hd__or2_2 _18865_ (.A(pcpi_rs2[15]),
    .B(_04605_),
    .X(_04609_));
 sky130_vsdinv _18866_ (.A(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__a21o_2 _18867_ (.A1(_11345_),
    .A2(_04605_),
    .B1(_04610_),
    .X(_02361_));
 sky130_vsdinv _18868_ (.A(_02362_),
    .Y(_04611_));
 sky130_fd_sc_hd__a22o_2 _18869_ (.A1(_11840_),
    .A2(_02362_),
    .B1(_12520_),
    .B2(_04611_),
    .X(_04612_));
 sky130_fd_sc_hd__o22a_2 _18870_ (.A1(_12516_),
    .A2(_04606_),
    .B1(_04607_),
    .B2(_04608_),
    .X(_04613_));
 sky130_fd_sc_hd__a2bb2oi_2 _18871_ (.A1_N(_04612_),
    .A2_N(_04613_),
    .B1(_04612_),
    .B2(_04613_),
    .Y(_02597_));
 sky130_fd_sc_hd__or2_2 _18872_ (.A(pcpi_rs2[16]),
    .B(_04609_),
    .X(_04614_));
 sky130_fd_sc_hd__o21ai_2 _18873_ (.A1(_02363_),
    .A2(_04610_),
    .B1(_04614_),
    .Y(_02364_));
 sky130_fd_sc_hd__o22ai_2 _18874_ (.A1(_12520_),
    .A2(_04611_),
    .B1(_04612_),
    .B2(_04613_),
    .Y(_04615_));
 sky130_fd_sc_hd__o2bb2a_2 _18875_ (.A1_N(pcpi_rs1[16]),
    .A2_N(_02365_),
    .B1(pcpi_rs1[16]),
    .B2(_02365_),
    .X(_04616_));
 sky130_fd_sc_hd__o2bb2a_2 _18876_ (.A1_N(_04615_),
    .A2_N(_04616_),
    .B1(_04615_),
    .B2(_04616_),
    .X(_02598_));
 sky130_fd_sc_hd__or2_2 _18877_ (.A(pcpi_rs2[17]),
    .B(_04614_),
    .X(_04617_));
 sky130_vsdinv _18878_ (.A(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__a21o_2 _18879_ (.A1(_11344_),
    .A2(_04614_),
    .B1(_04618_),
    .X(_02367_));
 sky130_fd_sc_hd__o2bb2a_2 _18880_ (.A1_N(_11837_),
    .A2_N(_02368_),
    .B1(_11837_),
    .B2(_02368_),
    .X(_04619_));
 sky130_fd_sc_hd__a22o_2 _18881_ (.A1(_11839_),
    .A2(_02365_),
    .B1(_04615_),
    .B2(_04616_),
    .X(_04620_));
 sky130_fd_sc_hd__a2bb2oi_2 _18882_ (.A1_N(_04619_),
    .A2_N(_04620_),
    .B1(_04619_),
    .B2(_04620_),
    .Y(_02599_));
 sky130_fd_sc_hd__or2_2 _18883_ (.A(pcpi_rs2[18]),
    .B(_04617_),
    .X(_04621_));
 sky130_fd_sc_hd__o21ai_2 _18884_ (.A1(_02369_),
    .A2(_04618_),
    .B1(_04621_),
    .Y(_02370_));
 sky130_vsdinv _18885_ (.A(_02371_),
    .Y(_04622_));
 sky130_fd_sc_hd__a22o_2 _18886_ (.A1(pcpi_rs1[18]),
    .A2(_02371_),
    .B1(_12534_),
    .B2(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__or2_2 _18887_ (.A(pcpi_rs1[17]),
    .B(_02368_),
    .X(_04624_));
 sky130_fd_sc_hd__a32o_2 _18888_ (.A1(pcpi_rs1[16]),
    .A2(_02365_),
    .A3(_04624_),
    .B1(_11838_),
    .B2(_02368_),
    .X(_04625_));
 sky130_fd_sc_hd__a31oi_2 _18889_ (.A1(_04616_),
    .A2(_04619_),
    .A3(_04615_),
    .B1(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__a2bb2oi_2 _18890_ (.A1_N(_04623_),
    .A2_N(_04626_),
    .B1(_04623_),
    .B2(_04626_),
    .Y(_02600_));
 sky130_fd_sc_hd__or2_2 _18891_ (.A(pcpi_rs2[19]),
    .B(_04621_),
    .X(_04627_));
 sky130_vsdinv _18892_ (.A(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__a21o_2 _18893_ (.A1(_11342_),
    .A2(_04621_),
    .B1(_04628_),
    .X(_02373_));
 sky130_vsdinv _18894_ (.A(_02374_),
    .Y(_04629_));
 sky130_fd_sc_hd__a22o_2 _18895_ (.A1(pcpi_rs1[19]),
    .A2(_02374_),
    .B1(_12541_),
    .B2(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__o22a_2 _18896_ (.A1(_12534_),
    .A2(_04622_),
    .B1(_04623_),
    .B2(_04626_),
    .X(_04631_));
 sky130_fd_sc_hd__a2bb2oi_2 _18897_ (.A1_N(_04630_),
    .A2_N(_04631_),
    .B1(_04630_),
    .B2(_04631_),
    .Y(_02601_));
 sky130_fd_sc_hd__or2_2 _18898_ (.A(pcpi_rs2[20]),
    .B(_04627_),
    .X(_04632_));
 sky130_fd_sc_hd__o21ai_2 _18899_ (.A1(_02375_),
    .A2(_04628_),
    .B1(_04632_),
    .Y(_02376_));
 sky130_vsdinv _18900_ (.A(_02377_),
    .Y(_04633_));
 sky130_fd_sc_hd__a22o_2 _18901_ (.A1(pcpi_rs1[20]),
    .A2(_02377_),
    .B1(_12545_),
    .B2(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__o22a_2 _18902_ (.A1(_12541_),
    .A2(_04629_),
    .B1(_04630_),
    .B2(_04631_),
    .X(_04635_));
 sky130_fd_sc_hd__a2bb2oi_2 _18903_ (.A1_N(_04634_),
    .A2_N(_04635_),
    .B1(_04634_),
    .B2(_04635_),
    .Y(_02603_));
 sky130_fd_sc_hd__or2_2 _18904_ (.A(pcpi_rs2[21]),
    .B(_04632_),
    .X(_04636_));
 sky130_vsdinv _18905_ (.A(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__a21o_2 _18906_ (.A1(_11340_),
    .A2(_04632_),
    .B1(_04637_),
    .X(_02379_));
 sky130_vsdinv _18907_ (.A(_02380_),
    .Y(_04638_));
 sky130_fd_sc_hd__a22o_2 _18908_ (.A1(pcpi_rs1[21]),
    .A2(_02380_),
    .B1(_12549_),
    .B2(_04638_),
    .X(_04639_));
 sky130_fd_sc_hd__o22a_2 _18909_ (.A1(_12545_),
    .A2(_04633_),
    .B1(_04634_),
    .B2(_04635_),
    .X(_04640_));
 sky130_fd_sc_hd__a2bb2oi_2 _18910_ (.A1_N(_04639_),
    .A2_N(_04640_),
    .B1(_04639_),
    .B2(_04640_),
    .Y(_02604_));
 sky130_fd_sc_hd__or2_2 _18911_ (.A(pcpi_rs2[22]),
    .B(_04636_),
    .X(_04641_));
 sky130_fd_sc_hd__o21ai_2 _18912_ (.A1(_02381_),
    .A2(_04637_),
    .B1(_04641_),
    .Y(_02382_));
 sky130_vsdinv _18913_ (.A(_02383_),
    .Y(_04642_));
 sky130_fd_sc_hd__a22o_2 _18914_ (.A1(pcpi_rs1[22]),
    .A2(_02383_),
    .B1(_12553_),
    .B2(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__o22a_2 _18915_ (.A1(_12549_),
    .A2(_04638_),
    .B1(_04639_),
    .B2(_04640_),
    .X(_04644_));
 sky130_fd_sc_hd__a2bb2oi_2 _18916_ (.A1_N(_04643_),
    .A2_N(_04644_),
    .B1(_04643_),
    .B2(_04644_),
    .Y(_02605_));
 sky130_fd_sc_hd__or2_2 _18917_ (.A(pcpi_rs2[23]),
    .B(_04641_),
    .X(_04645_));
 sky130_vsdinv _18918_ (.A(_04645_),
    .Y(_04646_));
 sky130_fd_sc_hd__a21o_2 _18919_ (.A1(_11339_),
    .A2(_04641_),
    .B1(_04646_),
    .X(_02385_));
 sky130_vsdinv _18920_ (.A(_02386_),
    .Y(_04647_));
 sky130_fd_sc_hd__a22o_2 _18921_ (.A1(pcpi_rs1[23]),
    .A2(_02386_),
    .B1(_12557_),
    .B2(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__o22a_2 _18922_ (.A1(_12553_),
    .A2(_04642_),
    .B1(_04643_),
    .B2(_04644_),
    .X(_04649_));
 sky130_fd_sc_hd__a2bb2oi_2 _18923_ (.A1_N(_04648_),
    .A2_N(_04649_),
    .B1(_04648_),
    .B2(_04649_),
    .Y(_02606_));
 sky130_fd_sc_hd__or2_2 _18924_ (.A(pcpi_rs2[24]),
    .B(_04645_),
    .X(_04650_));
 sky130_fd_sc_hd__o21ai_2 _18925_ (.A1(_02387_),
    .A2(_04646_),
    .B1(_04650_),
    .Y(_02388_));
 sky130_fd_sc_hd__o22ai_2 _18926_ (.A1(_12557_),
    .A2(_04647_),
    .B1(_04648_),
    .B2(_04649_),
    .Y(_04651_));
 sky130_fd_sc_hd__o2bb2a_2 _18927_ (.A1_N(_11827_),
    .A2_N(_02389_),
    .B1(_11827_),
    .B2(_02389_),
    .X(_04652_));
 sky130_fd_sc_hd__o2bb2a_2 _18928_ (.A1_N(_04651_),
    .A2_N(_04652_),
    .B1(_04651_),
    .B2(_04652_),
    .X(_02607_));
 sky130_fd_sc_hd__or2_2 _18929_ (.A(_11337_),
    .B(_04650_),
    .X(_04653_));
 sky130_vsdinv _18930_ (.A(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__a21o_2 _18931_ (.A1(_11337_),
    .A2(_04650_),
    .B1(_04654_),
    .X(_02391_));
 sky130_fd_sc_hd__o2bb2a_2 _18932_ (.A1_N(_11825_),
    .A2_N(_02392_),
    .B1(_11825_),
    .B2(_02392_),
    .X(_04655_));
 sky130_fd_sc_hd__a22o_2 _18933_ (.A1(_11828_),
    .A2(_02389_),
    .B1(_04651_),
    .B2(_04652_),
    .X(_04656_));
 sky130_fd_sc_hd__a2bb2oi_2 _18934_ (.A1_N(_04655_),
    .A2_N(_04656_),
    .B1(_04655_),
    .B2(_04656_),
    .Y(_02608_));
 sky130_fd_sc_hd__or2_2 _18935_ (.A(pcpi_rs2[26]),
    .B(_04653_),
    .X(_04657_));
 sky130_fd_sc_hd__o21ai_2 _18936_ (.A1(_02393_),
    .A2(_04654_),
    .B1(_04657_),
    .Y(_02394_));
 sky130_fd_sc_hd__or2_2 _18937_ (.A(_11824_),
    .B(_02392_),
    .X(_04658_));
 sky130_fd_sc_hd__a32o_2 _18938_ (.A1(_11827_),
    .A2(_02389_),
    .A3(_04658_),
    .B1(_11825_),
    .B2(_02392_),
    .X(_04659_));
 sky130_fd_sc_hd__a31o_2 _18939_ (.A1(_04652_),
    .A2(_04655_),
    .A3(_04651_),
    .B1(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__o2bb2a_2 _18940_ (.A1_N(_11821_),
    .A2_N(_02395_),
    .B1(_11821_),
    .B2(_02395_),
    .X(_04661_));
 sky130_fd_sc_hd__o2bb2a_2 _18941_ (.A1_N(_04660_),
    .A2_N(_04661_),
    .B1(_04660_),
    .B2(_04661_),
    .X(_02609_));
 sky130_fd_sc_hd__or2_2 _18942_ (.A(_11335_),
    .B(_04657_),
    .X(_04662_));
 sky130_vsdinv _18943_ (.A(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__a21o_2 _18944_ (.A1(_11335_),
    .A2(_04657_),
    .B1(_04663_),
    .X(_02397_));
 sky130_fd_sc_hd__o2bb2a_2 _18945_ (.A1_N(_11820_),
    .A2_N(_02398_),
    .B1(_11820_),
    .B2(_02398_),
    .X(_04664_));
 sky130_fd_sc_hd__a22o_2 _18946_ (.A1(_11822_),
    .A2(_02395_),
    .B1(_04660_),
    .B2(_04661_),
    .X(_04665_));
 sky130_fd_sc_hd__a2bb2oi_2 _18947_ (.A1_N(_04664_),
    .A2_N(_04665_),
    .B1(_04664_),
    .B2(_04665_),
    .Y(_02610_));
 sky130_fd_sc_hd__or2_2 _18948_ (.A(pcpi_rs2[28]),
    .B(_04662_),
    .X(_04666_));
 sky130_fd_sc_hd__o21ai_2 _18949_ (.A1(_02399_),
    .A2(_04663_),
    .B1(_04666_),
    .Y(_02400_));
 sky130_fd_sc_hd__or2_2 _18950_ (.A(_11819_),
    .B(_02398_),
    .X(_04667_));
 sky130_fd_sc_hd__a32o_2 _18951_ (.A1(_11822_),
    .A2(_02395_),
    .A3(_04667_),
    .B1(_11820_),
    .B2(_02398_),
    .X(_04668_));
 sky130_fd_sc_hd__a31o_2 _18952_ (.A1(_04661_),
    .A2(_04664_),
    .A3(_04660_),
    .B1(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__nor2_2 _18953_ (.A(pcpi_rs1[28]),
    .B(_02401_),
    .Y(_04670_));
 sky130_fd_sc_hd__a21oi_2 _18954_ (.A1(_11818_),
    .A2(_02401_),
    .B1(_04670_),
    .Y(_04671_));
 sky130_vsdinv _18955_ (.A(_04669_),
    .Y(_04672_));
 sky130_vsdinv _18956_ (.A(_04671_),
    .Y(_04673_));
 sky130_fd_sc_hd__o22a_2 _18957_ (.A1(_04669_),
    .A2(_04671_),
    .B1(_04672_),
    .B2(_04673_),
    .X(_02611_));
 sky130_fd_sc_hd__or2_2 _18958_ (.A(_11334_),
    .B(_04666_),
    .X(_04674_));
 sky130_vsdinv _18959_ (.A(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__a21o_2 _18960_ (.A1(_11334_),
    .A2(_04666_),
    .B1(_04675_),
    .X(_02403_));
 sky130_fd_sc_hd__o2bb2a_2 _18961_ (.A1_N(_11818_),
    .A2_N(_02401_),
    .B1(_04672_),
    .B2(_04670_),
    .X(_04676_));
 sky130_fd_sc_hd__nor2_2 _18962_ (.A(pcpi_rs1[29]),
    .B(_02404_),
    .Y(_04677_));
 sky130_fd_sc_hd__a21o_2 _18963_ (.A1(_11817_),
    .A2(_02404_),
    .B1(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__o2bb2a_2 _18964_ (.A1_N(_04676_),
    .A2_N(_04678_),
    .B1(_04676_),
    .B2(_04678_),
    .X(_02612_));
 sky130_fd_sc_hd__or2_2 _18965_ (.A(pcpi_rs2[30]),
    .B(_04674_),
    .X(_04679_));
 sky130_fd_sc_hd__o21ai_2 _18966_ (.A1(_02405_),
    .A2(_04675_),
    .B1(_04679_),
    .Y(_02406_));
 sky130_vsdinv _18967_ (.A(_02407_),
    .Y(_04680_));
 sky130_fd_sc_hd__a22o_2 _18968_ (.A1(_11816_),
    .A2(_02407_),
    .B1(_12595_),
    .B2(_04680_),
    .X(_04681_));
 sky130_fd_sc_hd__o2bb2a_2 _18969_ (.A1_N(_11817_),
    .A2_N(_02404_),
    .B1(_04676_),
    .B2(_04677_),
    .X(_04682_));
 sky130_fd_sc_hd__a2bb2oi_2 _18970_ (.A1_N(_04681_),
    .A2_N(_04682_),
    .B1(_04681_),
    .B2(_04682_),
    .Y(_02614_));
 sky130_fd_sc_hd__a32o_2 _18971_ (.A1(_02405_),
    .A2(_04675_),
    .A3(pcpi_rs2[31]),
    .B1(_10594_),
    .B2(_04679_),
    .X(_02408_));
 sky130_fd_sc_hd__o22ai_2 _18972_ (.A1(_12595_),
    .A2(_04680_),
    .B1(_04681_),
    .B2(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__a2bb2o_2 _18973_ (.A1_N(_10568_),
    .A2_N(_02409_),
    .B1(_10568_),
    .B2(_02409_),
    .X(_04684_));
 sky130_fd_sc_hd__a2bb2o_2 _18974_ (.A1_N(_04683_),
    .A2_N(_04684_),
    .B1(_04683_),
    .B2(_04684_),
    .X(_02615_));
 sky130_vsdinv _18975_ (.A(\pcpi_mul.rs1[1] ),
    .Y(_04685_));
 sky130_fd_sc_hd__buf_1 _18976_ (.A(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__buf_1 _18977_ (.A(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__buf_1 _18978_ (.A(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__buf_1 _18979_ (.A(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__buf_1 _18980_ (.A(_04689_),
    .X(_04690_));
 sky130_vsdinv _18981_ (.A(\pcpi_mul.rs2[1] ),
    .Y(_04691_));
 sky130_fd_sc_hd__buf_1 _18982_ (.A(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__buf_1 _18983_ (.A(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__buf_1 _18984_ (.A(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__buf_1 _18985_ (.A(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__o22a_2 _18986_ (.A1(_04539_),
    .A2(_04690_),
    .B1(_04695_),
    .B2(_04546_),
    .X(_04696_));
 sky130_fd_sc_hd__or4_2 _18987_ (.A(_04539_),
    .B(_04690_),
    .C(_04695_),
    .D(_04545_),
    .X(_04697_));
 sky130_fd_sc_hd__nor2b_2 _18988_ (.A(_04696_),
    .B_N(_04697_),
    .Y(_02624_));
 sky130_vsdinv _18989_ (.A(\pcpi_mul.rs1[2] ),
    .Y(_04698_));
 sky130_fd_sc_hd__buf_1 _18990_ (.A(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__buf_1 _18991_ (.A(_04699_),
    .X(_04700_));
 sky130_fd_sc_hd__buf_1 _18992_ (.A(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__buf_1 _18993_ (.A(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__buf_1 _18994_ (.A(_04688_),
    .X(_04703_));
 sky130_vsdinv _18995_ (.A(\pcpi_mul.rs2[2] ),
    .Y(_04704_));
 sky130_fd_sc_hd__buf_1 _18996_ (.A(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__buf_1 _18997_ (.A(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__buf_1 _18998_ (.A(_04542_),
    .X(_04707_));
 sky130_fd_sc_hd__o22a_2 _18999_ (.A1(_04693_),
    .A2(_04703_),
    .B1(_04706_),
    .B2(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__buf_1 _19000_ (.A(_04687_),
    .X(_04709_));
 sky130_fd_sc_hd__buf_1 _19001_ (.A(_04540_),
    .X(_04710_));
 sky130_fd_sc_hd__or4_2 _19002_ (.A(_04693_),
    .B(_04709_),
    .C(_04706_),
    .D(_04710_),
    .X(_04711_));
 sky130_vsdinv _19003_ (.A(_04711_),
    .Y(_04712_));
 sky130_fd_sc_hd__or2_2 _19004_ (.A(_04708_),
    .B(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__or3_2 _19005_ (.A(_04538_),
    .B(_04702_),
    .C(_04713_),
    .X(_04714_));
 sky130_vsdinv _19006_ (.A(_04714_),
    .Y(_04715_));
 sky130_fd_sc_hd__o21a_2 _19007_ (.A1(_04539_),
    .A2(_04702_),
    .B1(_04713_),
    .X(_04716_));
 sky130_fd_sc_hd__or2_2 _19008_ (.A(_04715_),
    .B(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__or2_2 _19009_ (.A(_04697_),
    .B(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__a21boi_2 _19010_ (.A1(_04697_),
    .A2(_04717_),
    .B1_N(_04718_),
    .Y(_02625_));
 sky130_fd_sc_hd__buf_1 _19011_ (.A(_04536_),
    .X(_04719_));
 sky130_vsdinv _19012_ (.A(\pcpi_mul.rs1[3] ),
    .Y(_04720_));
 sky130_fd_sc_hd__buf_1 _19013_ (.A(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__buf_1 _19014_ (.A(_04721_),
    .X(_04722_));
 sky130_fd_sc_hd__buf_1 _19015_ (.A(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__or2_2 _19016_ (.A(_04719_),
    .B(_04723_),
    .X(_04724_));
 sky130_fd_sc_hd__o22a_2 _19017_ (.A1(_04705_),
    .A2(_04687_),
    .B1(_04692_),
    .B2(_04700_),
    .X(_04725_));
 sky130_fd_sc_hd__and4_2 _19018_ (.A(_11635_),
    .B(_11954_),
    .C(_11641_),
    .D(_11951_),
    .X(_04726_));
 sky130_fd_sc_hd__nor2_2 _19019_ (.A(_04725_),
    .B(_04726_),
    .Y(_04727_));
 sky130_vsdinv _19020_ (.A(\pcpi_mul.rs2[3] ),
    .Y(_04728_));
 sky130_fd_sc_hd__buf_1 _19021_ (.A(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__buf_1 _19022_ (.A(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__nor2_2 _19023_ (.A(_04730_),
    .B(_04542_),
    .Y(_04731_));
 sky130_fd_sc_hd__a2bb2o_2 _19024_ (.A1_N(_04727_),
    .A2_N(_04731_),
    .B1(_04727_),
    .B2(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__or2_2 _19025_ (.A(_04724_),
    .B(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__a21bo_2 _19026_ (.A1(_04724_),
    .A2(_04732_),
    .B1_N(_04733_),
    .X(_04734_));
 sky130_vsdinv _19027_ (.A(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__o22a_2 _19028_ (.A1(_04715_),
    .A2(_04735_),
    .B1(_04714_),
    .B2(_04734_),
    .X(_04736_));
 sky130_fd_sc_hd__a2bb2o_2 _19029_ (.A1_N(_04712_),
    .A2_N(_04736_),
    .B1(_04712_),
    .B2(_04735_),
    .X(_04737_));
 sky130_fd_sc_hd__or2_2 _19030_ (.A(_04718_),
    .B(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__a21boi_2 _19031_ (.A1(_04718_),
    .A2(_04737_),
    .B1_N(_04738_),
    .Y(_02626_));
 sky130_vsdinv _19032_ (.A(\pcpi_mul.rs2[4] ),
    .Y(_04739_));
 sky130_fd_sc_hd__buf_1 _19033_ (.A(_04739_),
    .X(_04740_));
 sky130_vsdinv _19034_ (.A(\pcpi_mul.rs1[4] ),
    .Y(_04741_));
 sky130_fd_sc_hd__buf_1 _19035_ (.A(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__o22a_2 _19036_ (.A1(_04740_),
    .A2(_04541_),
    .B1(_04536_),
    .B2(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__buf_1 _19037_ (.A(_04535_),
    .X(_04744_));
 sky130_fd_sc_hd__buf_1 _19038_ (.A(_04741_),
    .X(_04745_));
 sky130_fd_sc_hd__or4_2 _19039_ (.A(_04740_),
    .B(_04541_),
    .C(_04744_),
    .D(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__or2b_2 _19040_ (.A(_04743_),
    .B_N(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__o22a_2 _19041_ (.A1(_04705_),
    .A2(_04699_),
    .B1(_04692_),
    .B2(_04721_),
    .X(_04748_));
 sky130_fd_sc_hd__and4_2 _19042_ (.A(_11634_),
    .B(_11950_),
    .C(_11640_),
    .D(_11947_),
    .X(_04749_));
 sky130_fd_sc_hd__nor2_2 _19043_ (.A(_04748_),
    .B(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__buf_1 _19044_ (.A(_04687_),
    .X(_04751_));
 sky130_fd_sc_hd__nor2_2 _19045_ (.A(_04729_),
    .B(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__a2bb2o_2 _19046_ (.A1_N(_04750_),
    .A2_N(_04752_),
    .B1(_04750_),
    .B2(_04752_),
    .X(_04753_));
 sky130_fd_sc_hd__or2_2 _19047_ (.A(_04747_),
    .B(_04753_),
    .X(_04754_));
 sky130_fd_sc_hd__a21bo_2 _19048_ (.A1(_04747_),
    .A2(_04753_),
    .B1_N(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__o2bb2a_2 _19049_ (.A1_N(_04733_),
    .A2_N(_04755_),
    .B1(_04733_),
    .B2(_04755_),
    .X(_04756_));
 sky130_vsdinv _19050_ (.A(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__a31o_2 _19051_ (.A1(\pcpi_mul.rs2[3] ),
    .A2(_11957_),
    .A3(_04727_),
    .B1(_04726_),
    .X(_04758_));
 sky130_vsdinv _19052_ (.A(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__a22o_2 _19053_ (.A1(_04757_),
    .A2(_04759_),
    .B1(_04756_),
    .B2(_04758_),
    .X(_04760_));
 sky130_fd_sc_hd__o22a_2 _19054_ (.A1(_04714_),
    .A2(_04734_),
    .B1(_04711_),
    .B2(_04734_),
    .X(_04761_));
 sky130_fd_sc_hd__or2_2 _19055_ (.A(_04760_),
    .B(_04761_),
    .X(_04762_));
 sky130_vsdinv _19056_ (.A(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__a21o_2 _19057_ (.A1(_04760_),
    .A2(_04761_),
    .B1(_04763_),
    .X(_04764_));
 sky130_fd_sc_hd__or2_2 _19058_ (.A(_04738_),
    .B(_04764_),
    .X(_04765_));
 sky130_vsdinv _19059_ (.A(_04765_),
    .Y(_04766_));
 sky130_fd_sc_hd__a21oi_2 _19060_ (.A1(_04738_),
    .A2(_04764_),
    .B1(_04766_),
    .Y(_02627_));
 sky130_fd_sc_hd__o22a_2 _19061_ (.A1(_04733_),
    .A2(_04755_),
    .B1(_04757_),
    .B2(_04759_),
    .X(_04767_));
 sky130_fd_sc_hd__a21oi_2 _19062_ (.A1(_04750_),
    .A2(_04752_),
    .B1(_04749_),
    .Y(_04768_));
 sky130_vsdinv _19063_ (.A(\pcpi_mul.rs1[5] ),
    .Y(_04769_));
 sky130_fd_sc_hd__buf_1 _19064_ (.A(_04769_),
    .X(_04770_));
 sky130_fd_sc_hd__or2_2 _19065_ (.A(_04744_),
    .B(_04770_),
    .X(_04771_));
 sky130_fd_sc_hd__and4_2 _19066_ (.A(_11630_),
    .B(_11953_),
    .C(_11626_),
    .D(_11956_),
    .X(_04772_));
 sky130_vsdinv _19067_ (.A(\pcpi_mul.rs2[5] ),
    .Y(_04773_));
 sky130_fd_sc_hd__buf_1 _19068_ (.A(_04773_),
    .X(_04774_));
 sky130_fd_sc_hd__o22a_2 _19069_ (.A1(_04740_),
    .A2(_04686_),
    .B1(_04774_),
    .B2(_04540_),
    .X(_04775_));
 sky130_fd_sc_hd__or2_2 _19070_ (.A(_04772_),
    .B(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__a2bb2o_2 _19071_ (.A1_N(_04771_),
    .A2_N(_04776_),
    .B1(_04771_),
    .B2(_04776_),
    .X(_04777_));
 sky130_fd_sc_hd__a2bb2o_2 _19072_ (.A1_N(_04746_),
    .A2_N(_04777_),
    .B1(_04746_),
    .B2(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__buf_1 _19073_ (.A(_04700_),
    .X(_04779_));
 sky130_fd_sc_hd__or2_2 _19074_ (.A(_04729_),
    .B(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__and4_2 _19075_ (.A(_11635_),
    .B(_11948_),
    .C(_11641_),
    .D(_11944_),
    .X(_04781_));
 sky130_fd_sc_hd__buf_1 _19076_ (.A(_04721_),
    .X(_04782_));
 sky130_fd_sc_hd__o22a_2 _19077_ (.A1(_04705_),
    .A2(_04782_),
    .B1(_04692_),
    .B2(_04742_),
    .X(_04783_));
 sky130_fd_sc_hd__or2_2 _19078_ (.A(_04781_),
    .B(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__a2bb2o_2 _19079_ (.A1_N(_04780_),
    .A2_N(_04784_),
    .B1(_04780_),
    .B2(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__a2bb2o_2 _19080_ (.A1_N(_04778_),
    .A2_N(_04785_),
    .B1(_04778_),
    .B2(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__a2bb2o_2 _19081_ (.A1_N(_04754_),
    .A2_N(_04786_),
    .B1(_04754_),
    .B2(_04786_),
    .X(_04787_));
 sky130_fd_sc_hd__a2bb2o_2 _19082_ (.A1_N(_04768_),
    .A2_N(_04787_),
    .B1(_04768_),
    .B2(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__or2_2 _19083_ (.A(_04767_),
    .B(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__a21bo_2 _19084_ (.A1(_04767_),
    .A2(_04788_),
    .B1_N(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__or2_2 _19085_ (.A(_04765_),
    .B(_04790_),
    .X(_04791_));
 sky130_vsdinv _19086_ (.A(\pcpi_mul.rs2[6] ),
    .Y(_04792_));
 sky130_fd_sc_hd__buf_1 _19087_ (.A(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__buf_1 _19088_ (.A(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__buf_1 _19089_ (.A(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__or2_2 _19090_ (.A(_04795_),
    .B(_04544_),
    .X(_04796_));
 sky130_fd_sc_hd__o21ba_2 _19091_ (.A1(_04780_),
    .A2(_04784_),
    .B1_N(_04781_),
    .X(_04797_));
 sky130_fd_sc_hd__and4_2 _19092_ (.A(_11634_),
    .B(_11944_),
    .C(_11640_),
    .D(_11941_),
    .X(_04798_));
 sky130_fd_sc_hd__o22a_2 _19093_ (.A1(_04705_),
    .A2(_04745_),
    .B1(_04691_),
    .B2(_04770_),
    .X(_04799_));
 sky130_fd_sc_hd__or2_2 _19094_ (.A(_04798_),
    .B(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__or2_2 _19095_ (.A(_04729_),
    .B(_04782_),
    .X(_04801_));
 sky130_fd_sc_hd__a2bb2o_2 _19096_ (.A1_N(_04800_),
    .A2_N(_04801_),
    .B1(_04800_),
    .B2(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__and4_2 _19097_ (.A(_11626_),
    .B(_11953_),
    .C(_11630_),
    .D(_11950_),
    .X(_04803_));
 sky130_fd_sc_hd__o22a_2 _19098_ (.A1(_04774_),
    .A2(_04685_),
    .B1(_04739_),
    .B2(_04699_),
    .X(_04804_));
 sky130_fd_sc_hd__or2_2 _19099_ (.A(_04803_),
    .B(_04804_),
    .X(_04805_));
 sky130_vsdinv _19100_ (.A(\pcpi_mul.rs1[6] ),
    .Y(_04806_));
 sky130_fd_sc_hd__buf_1 _19101_ (.A(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__or2_2 _19102_ (.A(_04744_),
    .B(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__a2bb2o_2 _19103_ (.A1_N(_04805_),
    .A2_N(_04808_),
    .B1(_04805_),
    .B2(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__o21ba_2 _19104_ (.A1(_04771_),
    .A2(_04776_),
    .B1_N(_04772_),
    .X(_04810_));
 sky130_fd_sc_hd__a2bb2o_2 _19105_ (.A1_N(_04809_),
    .A2_N(_04810_),
    .B1(_04809_),
    .B2(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__a2bb2o_2 _19106_ (.A1_N(_04802_),
    .A2_N(_04811_),
    .B1(_04802_),
    .B2(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__o22a_2 _19107_ (.A1(_04746_),
    .A2(_04777_),
    .B1(_04778_),
    .B2(_04785_),
    .X(_04813_));
 sky130_fd_sc_hd__a2bb2o_2 _19108_ (.A1_N(_04812_),
    .A2_N(_04813_),
    .B1(_04812_),
    .B2(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__a2bb2o_2 _19109_ (.A1_N(_04797_),
    .A2_N(_04814_),
    .B1(_04797_),
    .B2(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__or2_2 _19110_ (.A(_04796_),
    .B(_04815_),
    .X(_04816_));
 sky130_fd_sc_hd__a21bo_2 _19111_ (.A1(_04796_),
    .A2(_04815_),
    .B1_N(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__o22a_2 _19112_ (.A1(_04754_),
    .A2(_04786_),
    .B1(_04768_),
    .B2(_04787_),
    .X(_04818_));
 sky130_fd_sc_hd__or2_2 _19113_ (.A(_04817_),
    .B(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__a21bo_2 _19114_ (.A1(_04817_),
    .A2(_04818_),
    .B1_N(_04819_),
    .X(_04820_));
 sky130_fd_sc_hd__or2_2 _19115_ (.A(_04762_),
    .B(_04790_),
    .X(_04821_));
 sky130_fd_sc_hd__nand2_2 _19116_ (.A(_04789_),
    .B(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__a2bb2oi_2 _19117_ (.A1_N(_04820_),
    .A2_N(_04822_),
    .B1(_04820_),
    .B2(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__a2bb2oi_2 _19118_ (.A1_N(_04791_),
    .A2_N(_04823_),
    .B1(_04791_),
    .B2(_04823_),
    .Y(_02683_));
 sky130_fd_sc_hd__o22a_2 _19119_ (.A1(_04791_),
    .A2(_04823_),
    .B1(_04820_),
    .B2(_04821_),
    .X(_04824_));
 sky130_vsdinv _19120_ (.A(\pcpi_mul.rs2[7] ),
    .Y(_04825_));
 sky130_fd_sc_hd__buf_1 _19121_ (.A(_04825_),
    .X(_04826_));
 sky130_fd_sc_hd__buf_1 _19122_ (.A(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__buf_1 _19123_ (.A(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__buf_1 _19124_ (.A(_04793_),
    .X(_04829_));
 sky130_fd_sc_hd__buf_1 _19125_ (.A(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__o22a_2 _19126_ (.A1(_04828_),
    .A2(_04543_),
    .B1(_04830_),
    .B2(_04689_),
    .X(_04831_));
 sky130_fd_sc_hd__or4_2 _19127_ (.A(_04826_),
    .B(_04540_),
    .C(_04792_),
    .D(_04686_),
    .X(_04832_));
 sky130_fd_sc_hd__or2b_2 _19128_ (.A(_04831_),
    .B_N(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__o21ba_2 _19129_ (.A1(_04800_),
    .A2(_04801_),
    .B1_N(_04798_),
    .X(_04834_));
 sky130_fd_sc_hd__and4_2 _19130_ (.A(_11634_),
    .B(_11941_),
    .C(_11640_),
    .D(_11938_),
    .X(_04835_));
 sky130_fd_sc_hd__o22a_2 _19131_ (.A1(_04704_),
    .A2(_04770_),
    .B1(_04691_),
    .B2(_04807_),
    .X(_04836_));
 sky130_fd_sc_hd__or2_2 _19132_ (.A(_04835_),
    .B(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__or2_2 _19133_ (.A(_04729_),
    .B(_04742_),
    .X(_04838_));
 sky130_fd_sc_hd__a2bb2o_2 _19134_ (.A1_N(_04837_),
    .A2_N(_04838_),
    .B1(_04837_),
    .B2(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__and4_2 _19135_ (.A(\pcpi_mul.rs2[5] ),
    .B(\pcpi_mul.rs1[2] ),
    .C(\pcpi_mul.rs2[4] ),
    .D(\pcpi_mul.rs1[3] ),
    .X(_04840_));
 sky130_fd_sc_hd__o22a_2 _19136_ (.A1(_04773_),
    .A2(_04698_),
    .B1(_04739_),
    .B2(_04721_),
    .X(_04841_));
 sky130_fd_sc_hd__or2_2 _19137_ (.A(_04840_),
    .B(_04841_),
    .X(_04842_));
 sky130_vsdinv _19138_ (.A(\pcpi_mul.rs1[7] ),
    .Y(_04843_));
 sky130_fd_sc_hd__buf_1 _19139_ (.A(_04843_),
    .X(_04844_));
 sky130_fd_sc_hd__or2_2 _19140_ (.A(_04744_),
    .B(_04844_),
    .X(_04845_));
 sky130_fd_sc_hd__a2bb2o_2 _19141_ (.A1_N(_04842_),
    .A2_N(_04845_),
    .B1(_04842_),
    .B2(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__o21ba_2 _19142_ (.A1(_04805_),
    .A2(_04808_),
    .B1_N(_04803_),
    .X(_04847_));
 sky130_fd_sc_hd__a2bb2o_2 _19143_ (.A1_N(_04846_),
    .A2_N(_04847_),
    .B1(_04846_),
    .B2(_04847_),
    .X(_04848_));
 sky130_fd_sc_hd__a2bb2o_2 _19144_ (.A1_N(_04839_),
    .A2_N(_04848_),
    .B1(_04839_),
    .B2(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__o22a_2 _19145_ (.A1(_04809_),
    .A2(_04810_),
    .B1(_04802_),
    .B2(_04811_),
    .X(_04850_));
 sky130_fd_sc_hd__a2bb2o_2 _19146_ (.A1_N(_04849_),
    .A2_N(_04850_),
    .B1(_04849_),
    .B2(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__a2bb2o_2 _19147_ (.A1_N(_04834_),
    .A2_N(_04851_),
    .B1(_04834_),
    .B2(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__or2_2 _19148_ (.A(_04833_),
    .B(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__a21bo_2 _19149_ (.A1(_04833_),
    .A2(_04852_),
    .B1_N(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__or2_2 _19150_ (.A(_04816_),
    .B(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__a21bo_2 _19151_ (.A1(_04816_),
    .A2(_04854_),
    .B1_N(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__o22a_2 _19152_ (.A1(_04812_),
    .A2(_04813_),
    .B1(_04797_),
    .B2(_04814_),
    .X(_04857_));
 sky130_fd_sc_hd__or2_2 _19153_ (.A(_04856_),
    .B(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__a21bo_2 _19154_ (.A1(_04856_),
    .A2(_04857_),
    .B1_N(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__or2_2 _19155_ (.A(_04789_),
    .B(_04820_),
    .X(_04860_));
 sky130_fd_sc_hd__nand2_2 _19156_ (.A(_04819_),
    .B(_04860_),
    .Y(_04861_));
 sky130_fd_sc_hd__a2bb2oi_2 _19157_ (.A1_N(_04859_),
    .A2_N(_04861_),
    .B1(_04859_),
    .B2(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__a2bb2oi_2 _19158_ (.A1_N(_04824_),
    .A2_N(_04862_),
    .B1(_04824_),
    .B2(_04862_),
    .Y(_02684_));
 sky130_fd_sc_hd__o22a_2 _19159_ (.A1(_04824_),
    .A2(_04862_),
    .B1(_04859_),
    .B2(_04860_),
    .X(_04863_));
 sky130_fd_sc_hd__and4_2 _19160_ (.A(_11622_),
    .B(\pcpi_mul.rs1[1] ),
    .C(\pcpi_mul.rs2[8] ),
    .D(\pcpi_mul.rs1[0] ),
    .X(_04864_));
 sky130_vsdinv _19161_ (.A(\pcpi_mul.rs2[8] ),
    .Y(_04865_));
 sky130_fd_sc_hd__o22a_2 _19162_ (.A1(_04825_),
    .A2(_04685_),
    .B1(_04865_),
    .B2(_04540_),
    .X(_04866_));
 sky130_fd_sc_hd__or2_2 _19163_ (.A(_04864_),
    .B(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__or2_2 _19164_ (.A(_04792_),
    .B(_04698_),
    .X(_04868_));
 sky130_fd_sc_hd__a2bb2o_2 _19165_ (.A1_N(_04867_),
    .A2_N(_04868_),
    .B1(_04867_),
    .B2(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__or2_2 _19166_ (.A(_04832_),
    .B(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__a21bo_2 _19167_ (.A1(_04832_),
    .A2(_04869_),
    .B1_N(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__o21ba_2 _19168_ (.A1(_04837_),
    .A2(_04838_),
    .B1_N(_04835_),
    .X(_04872_));
 sky130_fd_sc_hd__and4_2 _19169_ (.A(_11634_),
    .B(\pcpi_mul.rs1[6] ),
    .C(_11640_),
    .D(\pcpi_mul.rs1[7] ),
    .X(_04873_));
 sky130_fd_sc_hd__o22a_2 _19170_ (.A1(_04704_),
    .A2(_04806_),
    .B1(_04691_),
    .B2(_04843_),
    .X(_04874_));
 sky130_fd_sc_hd__or2_2 _19171_ (.A(_04873_),
    .B(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__buf_1 _19172_ (.A(_04770_),
    .X(_04876_));
 sky130_fd_sc_hd__or2_2 _19173_ (.A(_04728_),
    .B(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__a2bb2o_2 _19174_ (.A1_N(_04875_),
    .A2_N(_04877_),
    .B1(_04875_),
    .B2(_04877_),
    .X(_04878_));
 sky130_vsdinv _19175_ (.A(\pcpi_mul.rs1[8] ),
    .Y(_04879_));
 sky130_fd_sc_hd__or2_2 _19176_ (.A(_04535_),
    .B(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__and4_2 _19177_ (.A(\pcpi_mul.rs2[4] ),
    .B(\pcpi_mul.rs1[4] ),
    .C(\pcpi_mul.rs2[5] ),
    .D(\pcpi_mul.rs1[3] ),
    .X(_04881_));
 sky130_fd_sc_hd__o22a_2 _19178_ (.A1(_04739_),
    .A2(_04741_),
    .B1(_04774_),
    .B2(_04720_),
    .X(_04882_));
 sky130_fd_sc_hd__or2_2 _19179_ (.A(_04881_),
    .B(_04882_),
    .X(_04883_));
 sky130_fd_sc_hd__a2bb2o_2 _19180_ (.A1_N(_04880_),
    .A2_N(_04883_),
    .B1(_04880_),
    .B2(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__o21ba_2 _19181_ (.A1(_04842_),
    .A2(_04845_),
    .B1_N(_04840_),
    .X(_04885_));
 sky130_fd_sc_hd__a2bb2o_2 _19182_ (.A1_N(_04884_),
    .A2_N(_04885_),
    .B1(_04884_),
    .B2(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__a2bb2o_2 _19183_ (.A1_N(_04878_),
    .A2_N(_04886_),
    .B1(_04878_),
    .B2(_04886_),
    .X(_04887_));
 sky130_fd_sc_hd__o22a_2 _19184_ (.A1(_04846_),
    .A2(_04847_),
    .B1(_04839_),
    .B2(_04848_),
    .X(_04888_));
 sky130_fd_sc_hd__a2bb2o_2 _19185_ (.A1_N(_04887_),
    .A2_N(_04888_),
    .B1(_04887_),
    .B2(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__a2bb2o_2 _19186_ (.A1_N(_04872_),
    .A2_N(_04889_),
    .B1(_04872_),
    .B2(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__nor2_2 _19187_ (.A(_04871_),
    .B(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__a21o_2 _19188_ (.A1(_04871_),
    .A2(_04890_),
    .B1(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__or2_2 _19189_ (.A(_04853_),
    .B(_04892_),
    .X(_04893_));
 sky130_fd_sc_hd__a21bo_2 _19190_ (.A1(_04853_),
    .A2(_04892_),
    .B1_N(_04893_),
    .X(_04894_));
 sky130_fd_sc_hd__o22a_2 _19191_ (.A1(_04849_),
    .A2(_04850_),
    .B1(_04834_),
    .B2(_04851_),
    .X(_04895_));
 sky130_fd_sc_hd__a2bb2o_2 _19192_ (.A1_N(_04855_),
    .A2_N(_04895_),
    .B1(_04855_),
    .B2(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__a2bb2o_2 _19193_ (.A1_N(_04894_),
    .A2_N(_04896_),
    .B1(_04894_),
    .B2(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__o21ai_2 _19194_ (.A1(_04819_),
    .A2(_04859_),
    .B1(_04858_),
    .Y(_04898_));
 sky130_fd_sc_hd__a2bb2oi_2 _19195_ (.A1_N(_04897_),
    .A2_N(_04898_),
    .B1(_04897_),
    .B2(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__a2bb2oi_2 _19196_ (.A1_N(_04863_),
    .A2_N(_04899_),
    .B1(_04863_),
    .B2(_04899_),
    .Y(_02685_));
 sky130_fd_sc_hd__or2_2 _19197_ (.A(_04858_),
    .B(_04897_),
    .X(_04900_));
 sky130_vsdinv _19198_ (.A(\pcpi_mul.rs2[9] ),
    .Y(_04901_));
 sky130_fd_sc_hd__buf_1 _19199_ (.A(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__buf_1 _19200_ (.A(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__or2_2 _19201_ (.A(_04903_),
    .B(_04546_),
    .X(_04904_));
 sky130_fd_sc_hd__and4_2 _19202_ (.A(\pcpi_mul.rs2[8] ),
    .B(_11953_),
    .C(\pcpi_mul.rs2[7] ),
    .D(\pcpi_mul.rs1[2] ),
    .X(_04905_));
 sky130_fd_sc_hd__o22a_2 _19203_ (.A1(_04865_),
    .A2(_04685_),
    .B1(_04825_),
    .B2(_04698_),
    .X(_04906_));
 sky130_fd_sc_hd__or2_2 _19204_ (.A(_04905_),
    .B(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__or2_2 _19205_ (.A(_04792_),
    .B(_04720_),
    .X(_04908_));
 sky130_fd_sc_hd__a2bb2o_2 _19206_ (.A1_N(_04907_),
    .A2_N(_04908_),
    .B1(_04907_),
    .B2(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__o21ba_2 _19207_ (.A1(_04867_),
    .A2(_04868_),
    .B1_N(_04864_),
    .X(_04910_));
 sky130_fd_sc_hd__or2_2 _19208_ (.A(_04909_),
    .B(_04910_),
    .X(_04911_));
 sky130_vsdinv _19209_ (.A(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__a21o_2 _19210_ (.A1(_04909_),
    .A2(_04910_),
    .B1(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__or2_2 _19211_ (.A(_04870_),
    .B(_04913_),
    .X(_04914_));
 sky130_vsdinv _19212_ (.A(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__a21o_2 _19213_ (.A1(_04870_),
    .A2(_04913_),
    .B1(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__o21ba_2 _19214_ (.A1(_04875_),
    .A2(_04877_),
    .B1_N(_04873_),
    .X(_04917_));
 sky130_fd_sc_hd__and4_2 _19215_ (.A(_11634_),
    .B(\pcpi_mul.rs1[7] ),
    .C(_11640_),
    .D(\pcpi_mul.rs1[8] ),
    .X(_04918_));
 sky130_fd_sc_hd__o22a_2 _19216_ (.A1(_04704_),
    .A2(_04843_),
    .B1(_04691_),
    .B2(_04879_),
    .X(_04919_));
 sky130_fd_sc_hd__or2_2 _19217_ (.A(_04918_),
    .B(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__or2_2 _19218_ (.A(_04728_),
    .B(_04807_),
    .X(_04921_));
 sky130_fd_sc_hd__a2bb2o_2 _19219_ (.A1_N(_04920_),
    .A2_N(_04921_),
    .B1(_04920_),
    .B2(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__and4_2 _19220_ (.A(\pcpi_mul.rs2[5] ),
    .B(\pcpi_mul.rs1[4] ),
    .C(\pcpi_mul.rs2[4] ),
    .D(\pcpi_mul.rs1[5] ),
    .X(_04923_));
 sky130_fd_sc_hd__o22a_2 _19221_ (.A1(_04773_),
    .A2(_04741_),
    .B1(_04739_),
    .B2(_04769_),
    .X(_04924_));
 sky130_fd_sc_hd__or2_2 _19222_ (.A(_04923_),
    .B(_04924_),
    .X(_04925_));
 sky130_vsdinv _19223_ (.A(\pcpi_mul.rs1[9] ),
    .Y(_04926_));
 sky130_fd_sc_hd__or2_2 _19224_ (.A(_04744_),
    .B(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__a2bb2o_2 _19225_ (.A1_N(_04925_),
    .A2_N(_04927_),
    .B1(_04925_),
    .B2(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__o21ba_2 _19226_ (.A1(_04880_),
    .A2(_04883_),
    .B1_N(_04881_),
    .X(_04929_));
 sky130_fd_sc_hd__a2bb2o_2 _19227_ (.A1_N(_04928_),
    .A2_N(_04929_),
    .B1(_04928_),
    .B2(_04929_),
    .X(_04930_));
 sky130_fd_sc_hd__a2bb2o_2 _19228_ (.A1_N(_04922_),
    .A2_N(_04930_),
    .B1(_04922_),
    .B2(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__o22a_2 _19229_ (.A1(_04884_),
    .A2(_04885_),
    .B1(_04878_),
    .B2(_04886_),
    .X(_04932_));
 sky130_fd_sc_hd__a2bb2o_2 _19230_ (.A1_N(_04931_),
    .A2_N(_04932_),
    .B1(_04931_),
    .B2(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__a2bb2o_2 _19231_ (.A1_N(_04917_),
    .A2_N(_04933_),
    .B1(_04917_),
    .B2(_04933_),
    .X(_04934_));
 sky130_fd_sc_hd__or2_2 _19232_ (.A(_04916_),
    .B(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__a21boi_2 _19233_ (.A1(_04916_),
    .A2(_04934_),
    .B1_N(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__nand2_2 _19234_ (.A(_04891_),
    .B(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__o21ai_2 _19235_ (.A1(_04891_),
    .A2(_04936_),
    .B1(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__or2_2 _19236_ (.A(_04904_),
    .B(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__a21bo_2 _19237_ (.A1(_04904_),
    .A2(_04938_),
    .B1_N(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__o22a_2 _19238_ (.A1(_04887_),
    .A2(_04888_),
    .B1(_04872_),
    .B2(_04889_),
    .X(_04941_));
 sky130_fd_sc_hd__a2bb2o_2 _19239_ (.A1_N(_04893_),
    .A2_N(_04941_),
    .B1(_04893_),
    .B2(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__a2bb2o_2 _19240_ (.A1_N(_04940_),
    .A2_N(_04942_),
    .B1(_04940_),
    .B2(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__o22a_2 _19241_ (.A1(_04855_),
    .A2(_04895_),
    .B1(_04894_),
    .B2(_04896_),
    .X(_04944_));
 sky130_fd_sc_hd__or2_2 _19242_ (.A(_04943_),
    .B(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__a21bo_2 _19243_ (.A1(_04943_),
    .A2(_04944_),
    .B1_N(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__a2bb2o_2 _19244_ (.A1_N(_04900_),
    .A2_N(_04946_),
    .B1(_04900_),
    .B2(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__o32a_2 _19245_ (.A1(_04819_),
    .A2(_04859_),
    .A3(_04897_),
    .B1(_04863_),
    .B2(_04899_),
    .X(_04948_));
 sky130_fd_sc_hd__a2bb2oi_2 _19246_ (.A1_N(_04947_),
    .A2_N(_04948_),
    .B1(_04947_),
    .B2(_04948_),
    .Y(_02686_));
 sky130_vsdinv _19247_ (.A(\pcpi_mul.rs2[10] ),
    .Y(_04949_));
 sky130_fd_sc_hd__buf_1 _19248_ (.A(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__buf_1 _19249_ (.A(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__o22a_2 _19250_ (.A1(_04951_),
    .A2(_04545_),
    .B1(_04903_),
    .B2(_04690_),
    .X(_04952_));
 sky130_fd_sc_hd__buf_1 _19251_ (.A(_04901_),
    .X(_04953_));
 sky130_fd_sc_hd__or4_2 _19252_ (.A(_04950_),
    .B(_04542_),
    .C(_04953_),
    .D(_04688_),
    .X(_04954_));
 sky130_fd_sc_hd__or2b_2 _19253_ (.A(_04952_),
    .B_N(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__o21ba_2 _19254_ (.A1(_04920_),
    .A2(_04921_),
    .B1_N(_04918_),
    .X(_04956_));
 sky130_fd_sc_hd__and4_2 _19255_ (.A(_11635_),
    .B(\pcpi_mul.rs1[8] ),
    .C(_11641_),
    .D(\pcpi_mul.rs1[9] ),
    .X(_04957_));
 sky130_fd_sc_hd__buf_1 _19256_ (.A(_04879_),
    .X(_04958_));
 sky130_fd_sc_hd__o22a_2 _19257_ (.A1(_04705_),
    .A2(_04958_),
    .B1(_04692_),
    .B2(_04926_),
    .X(_04959_));
 sky130_fd_sc_hd__or2_2 _19258_ (.A(_04957_),
    .B(_04959_),
    .X(_04960_));
 sky130_fd_sc_hd__or2_2 _19259_ (.A(_04729_),
    .B(_04844_),
    .X(_04961_));
 sky130_fd_sc_hd__a2bb2o_2 _19260_ (.A1_N(_04960_),
    .A2_N(_04961_),
    .B1(_04960_),
    .B2(_04961_),
    .X(_04962_));
 sky130_vsdinv _19261_ (.A(\pcpi_mul.rs1[10] ),
    .Y(_04963_));
 sky130_fd_sc_hd__or2_2 _19262_ (.A(_04744_),
    .B(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__and4_2 _19263_ (.A(_11626_),
    .B(\pcpi_mul.rs1[5] ),
    .C(_11630_),
    .D(\pcpi_mul.rs1[6] ),
    .X(_04965_));
 sky130_fd_sc_hd__o22a_2 _19264_ (.A1(_04774_),
    .A2(_04769_),
    .B1(_04740_),
    .B2(_04806_),
    .X(_04966_));
 sky130_fd_sc_hd__or2_2 _19265_ (.A(_04965_),
    .B(_04966_),
    .X(_04967_));
 sky130_fd_sc_hd__a2bb2o_2 _19266_ (.A1_N(_04964_),
    .A2_N(_04967_),
    .B1(_04964_),
    .B2(_04967_),
    .X(_04968_));
 sky130_fd_sc_hd__o21ba_2 _19267_ (.A1(_04925_),
    .A2(_04927_),
    .B1_N(_04923_),
    .X(_04969_));
 sky130_fd_sc_hd__a2bb2o_2 _19268_ (.A1_N(_04968_),
    .A2_N(_04969_),
    .B1(_04968_),
    .B2(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__a2bb2o_2 _19269_ (.A1_N(_04962_),
    .A2_N(_04970_),
    .B1(_04962_),
    .B2(_04970_),
    .X(_04971_));
 sky130_fd_sc_hd__o22a_2 _19270_ (.A1(_04928_),
    .A2(_04929_),
    .B1(_04922_),
    .B2(_04930_),
    .X(_04972_));
 sky130_fd_sc_hd__a2bb2o_2 _19271_ (.A1_N(_04971_),
    .A2_N(_04972_),
    .B1(_04971_),
    .B2(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__a2bb2o_2 _19272_ (.A1_N(_04956_),
    .A2_N(_04973_),
    .B1(_04956_),
    .B2(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__buf_1 _19273_ (.A(_04745_),
    .X(_04975_));
 sky130_fd_sc_hd__or2_2 _19274_ (.A(_04793_),
    .B(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__buf_1 _19275_ (.A(_04865_),
    .X(_04977_));
 sky130_fd_sc_hd__o22a_2 _19276_ (.A1(_04977_),
    .A2(_04699_),
    .B1(_04826_),
    .B2(_04721_),
    .X(_04978_));
 sky130_fd_sc_hd__and4_2 _19277_ (.A(_11618_),
    .B(_11950_),
    .C(_11622_),
    .D(_11947_),
    .X(_04979_));
 sky130_fd_sc_hd__or2_2 _19278_ (.A(_04978_),
    .B(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__a2bb2o_2 _19279_ (.A1_N(_04976_),
    .A2_N(_04980_),
    .B1(_04976_),
    .B2(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__o21ba_2 _19280_ (.A1(_04907_),
    .A2(_04908_),
    .B1_N(_04905_),
    .X(_04982_));
 sky130_fd_sc_hd__or2_2 _19281_ (.A(_04981_),
    .B(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__a21bo_2 _19282_ (.A1(_04981_),
    .A2(_04982_),
    .B1_N(_04983_),
    .X(_04984_));
 sky130_fd_sc_hd__or2_2 _19283_ (.A(_04912_),
    .B(_04915_),
    .X(_04985_));
 sky130_fd_sc_hd__a2bb2oi_2 _19284_ (.A1_N(_04984_),
    .A2_N(_04985_),
    .B1(_04984_),
    .B2(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__a2bb2o_2 _19285_ (.A1_N(_04974_),
    .A2_N(_04986_),
    .B1(_04974_),
    .B2(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__or2_2 _19286_ (.A(_04935_),
    .B(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__a21bo_2 _19287_ (.A1(_04935_),
    .A2(_04987_),
    .B1_N(_04988_),
    .X(_04989_));
 sky130_fd_sc_hd__or2_2 _19288_ (.A(_04955_),
    .B(_04989_),
    .X(_04990_));
 sky130_fd_sc_hd__a21bo_2 _19289_ (.A1(_04955_),
    .A2(_04989_),
    .B1_N(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__a2bb2o_2 _19290_ (.A1_N(_04939_),
    .A2_N(_04991_),
    .B1(_04939_),
    .B2(_04991_),
    .X(_04992_));
 sky130_fd_sc_hd__o22a_2 _19291_ (.A1(_04931_),
    .A2(_04932_),
    .B1(_04917_),
    .B2(_04933_),
    .X(_04993_));
 sky130_fd_sc_hd__or2_2 _19292_ (.A(_04937_),
    .B(_04993_),
    .X(_04994_));
 sky130_fd_sc_hd__a21bo_2 _19293_ (.A1(_04937_),
    .A2(_04993_),
    .B1_N(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__a2bb2o_2 _19294_ (.A1_N(_04992_),
    .A2_N(_04995_),
    .B1(_04992_),
    .B2(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__o22a_2 _19295_ (.A1(_04893_),
    .A2(_04941_),
    .B1(_04940_),
    .B2(_04942_),
    .X(_04997_));
 sky130_fd_sc_hd__or2_2 _19296_ (.A(_04996_),
    .B(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__a21bo_2 _19297_ (.A1(_04996_),
    .A2(_04997_),
    .B1_N(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__a2bb2o_2 _19298_ (.A1_N(_04945_),
    .A2_N(_04999_),
    .B1(_04945_),
    .B2(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__o22a_2 _19299_ (.A1(_04900_),
    .A2(_04946_),
    .B1(_04947_),
    .B2(_04948_),
    .X(_05001_));
 sky130_fd_sc_hd__a2bb2oi_2 _19300_ (.A1_N(_05000_),
    .A2_N(_05001_),
    .B1(_05000_),
    .B2(_05001_),
    .Y(_02629_));
 sky130_fd_sc_hd__o22a_2 _19301_ (.A1(_04971_),
    .A2(_04972_),
    .B1(_04956_),
    .B2(_04973_),
    .X(_05002_));
 sky130_fd_sc_hd__or2_2 _19302_ (.A(_04988_),
    .B(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__a21bo_2 _19303_ (.A1(_04988_),
    .A2(_05002_),
    .B1_N(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__or2_2 _19304_ (.A(_04901_),
    .B(_04779_),
    .X(_05005_));
 sky130_fd_sc_hd__and4_2 _19305_ (.A(\pcpi_mul.rs2[10] ),
    .B(_11954_),
    .C(\pcpi_mul.rs2[11] ),
    .D(_11956_),
    .X(_05006_));
 sky130_vsdinv _19306_ (.A(\pcpi_mul.rs2[11] ),
    .Y(_05007_));
 sky130_fd_sc_hd__o22a_2 _19307_ (.A1(_04949_),
    .A2(_04686_),
    .B1(_05007_),
    .B2(_04541_),
    .X(_05008_));
 sky130_fd_sc_hd__or2_2 _19308_ (.A(_05006_),
    .B(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__a2bb2o_2 _19309_ (.A1_N(_05005_),
    .A2_N(_05009_),
    .B1(_05005_),
    .B2(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__o21ba_2 _19310_ (.A1(_04960_),
    .A2(_04961_),
    .B1_N(_04957_),
    .X(_05011_));
 sky130_fd_sc_hd__and4_2 _19311_ (.A(_11635_),
    .B(_11930_),
    .C(_11641_),
    .D(\pcpi_mul.rs1[10] ),
    .X(_05012_));
 sky130_fd_sc_hd__buf_1 _19312_ (.A(_04926_),
    .X(_05013_));
 sky130_fd_sc_hd__buf_1 _19313_ (.A(_04963_),
    .X(_05014_));
 sky130_fd_sc_hd__o22a_2 _19314_ (.A1(_04706_),
    .A2(_05013_),
    .B1(_04692_),
    .B2(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__or2_2 _19315_ (.A(_05012_),
    .B(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__buf_1 _19316_ (.A(_04958_),
    .X(_05017_));
 sky130_fd_sc_hd__or2_2 _19317_ (.A(_04730_),
    .B(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__a2bb2o_2 _19318_ (.A1_N(_05016_),
    .A2_N(_05018_),
    .B1(_05016_),
    .B2(_05018_),
    .X(_05019_));
 sky130_vsdinv _19319_ (.A(\pcpi_mul.rs1[11] ),
    .Y(_05020_));
 sky130_fd_sc_hd__or2_2 _19320_ (.A(_04536_),
    .B(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__and4_2 _19321_ (.A(_11626_),
    .B(_11938_),
    .C(_11630_),
    .D(_11936_),
    .X(_05022_));
 sky130_fd_sc_hd__o22a_2 _19322_ (.A1(_04774_),
    .A2(_04807_),
    .B1(_04740_),
    .B2(_04844_),
    .X(_05023_));
 sky130_fd_sc_hd__or2_2 _19323_ (.A(_05022_),
    .B(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__a2bb2o_2 _19324_ (.A1_N(_05021_),
    .A2_N(_05024_),
    .B1(_05021_),
    .B2(_05024_),
    .X(_05025_));
 sky130_fd_sc_hd__o21ba_2 _19325_ (.A1(_04964_),
    .A2(_04967_),
    .B1_N(_04965_),
    .X(_05026_));
 sky130_fd_sc_hd__a2bb2o_2 _19326_ (.A1_N(_05025_),
    .A2_N(_05026_),
    .B1(_05025_),
    .B2(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__a2bb2o_2 _19327_ (.A1_N(_05019_),
    .A2_N(_05027_),
    .B1(_05019_),
    .B2(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__o22a_2 _19328_ (.A1(_04968_),
    .A2(_04969_),
    .B1(_04962_),
    .B2(_04970_),
    .X(_05029_));
 sky130_fd_sc_hd__a2bb2o_2 _19329_ (.A1_N(_05028_),
    .A2_N(_05029_),
    .B1(_05028_),
    .B2(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__a2bb2o_2 _19330_ (.A1_N(_05011_),
    .A2_N(_05030_),
    .B1(_05011_),
    .B2(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__o21ba_2 _19331_ (.A1(_04976_),
    .A2(_04980_),
    .B1_N(_04979_),
    .X(_05032_));
 sky130_fd_sc_hd__or2_2 _19332_ (.A(_04793_),
    .B(_04876_),
    .X(_05033_));
 sky130_fd_sc_hd__o22a_2 _19333_ (.A1(_04977_),
    .A2(_04782_),
    .B1(_04826_),
    .B2(_04745_),
    .X(_05034_));
 sky130_fd_sc_hd__and4_2 _19334_ (.A(_11618_),
    .B(_11947_),
    .C(_11622_),
    .D(_11944_),
    .X(_05035_));
 sky130_fd_sc_hd__or2_2 _19335_ (.A(_05034_),
    .B(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__a2bb2o_2 _19336_ (.A1_N(_05033_),
    .A2_N(_05036_),
    .B1(_05033_),
    .B2(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__a2bb2o_2 _19337_ (.A1_N(_04954_),
    .A2_N(_05037_),
    .B1(_04954_),
    .B2(_05037_),
    .X(_05038_));
 sky130_fd_sc_hd__a2bb2o_2 _19338_ (.A1_N(_05032_),
    .A2_N(_05038_),
    .B1(_05032_),
    .B2(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__o21ai_2 _19339_ (.A1(_04911_),
    .A2(_04984_),
    .B1(_04983_),
    .Y(_05040_));
 sky130_fd_sc_hd__a2bb2oi_2 _19340_ (.A1_N(_05039_),
    .A2_N(_05040_),
    .B1(_05039_),
    .B2(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__a2bb2o_2 _19341_ (.A1_N(_05031_),
    .A2_N(_05041_),
    .B1(_05031_),
    .B2(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__o22a_2 _19342_ (.A1(_04974_),
    .A2(_04986_),
    .B1(_04914_),
    .B2(_04984_),
    .X(_05043_));
 sky130_fd_sc_hd__or2_2 _19343_ (.A(_05042_),
    .B(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__a21bo_2 _19344_ (.A1(_05042_),
    .A2(_05043_),
    .B1_N(_05044_),
    .X(_05045_));
 sky130_fd_sc_hd__or2_2 _19345_ (.A(_05010_),
    .B(_05045_),
    .X(_05046_));
 sky130_fd_sc_hd__a21bo_2 _19346_ (.A1(_05010_),
    .A2(_05045_),
    .B1_N(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__a2bb2o_2 _19347_ (.A1_N(_04990_),
    .A2_N(_05047_),
    .B1(_04990_),
    .B2(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__a2bb2o_2 _19348_ (.A1_N(_05004_),
    .A2_N(_05048_),
    .B1(_05004_),
    .B2(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__o22a_2 _19349_ (.A1(_04939_),
    .A2(_04991_),
    .B1(_04992_),
    .B2(_04995_),
    .X(_05050_));
 sky130_fd_sc_hd__a2bb2o_2 _19350_ (.A1_N(_05049_),
    .A2_N(_05050_),
    .B1(_05049_),
    .B2(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__a2bb2o_2 _19351_ (.A1_N(_04994_),
    .A2_N(_05051_),
    .B1(_04994_),
    .B2(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__a2bb2o_2 _19352_ (.A1_N(_04998_),
    .A2_N(_05052_),
    .B1(_04998_),
    .B2(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__o22a_2 _19353_ (.A1(_04945_),
    .A2(_04999_),
    .B1(_05000_),
    .B2(_05001_),
    .X(_05054_));
 sky130_fd_sc_hd__a2bb2oi_2 _19354_ (.A1_N(_05053_),
    .A2_N(_05054_),
    .B1(_05053_),
    .B2(_05054_),
    .Y(_02630_));
 sky130_vsdinv _19355_ (.A(\pcpi_mul.rs2[12] ),
    .Y(_05055_));
 sky130_fd_sc_hd__buf_1 _19356_ (.A(_05055_),
    .X(_05056_));
 sky130_fd_sc_hd__buf_1 _19357_ (.A(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__or2_2 _19358_ (.A(_05057_),
    .B(_04544_),
    .X(_05058_));
 sky130_fd_sc_hd__or2_2 _19359_ (.A(_04902_),
    .B(_04723_),
    .X(_05059_));
 sky130_fd_sc_hd__buf_1 _19360_ (.A(_05007_),
    .X(_05060_));
 sky130_fd_sc_hd__buf_1 _19361_ (.A(_04700_),
    .X(_05061_));
 sky130_fd_sc_hd__o22a_2 _19362_ (.A1(_05060_),
    .A2(_04688_),
    .B1(_04950_),
    .B2(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__and4_2 _19363_ (.A(_11613_),
    .B(_11955_),
    .C(_11616_),
    .D(_11952_),
    .X(_05063_));
 sky130_fd_sc_hd__or2_2 _19364_ (.A(_05062_),
    .B(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__a2bb2o_2 _19365_ (.A1_N(_05059_),
    .A2_N(_05064_),
    .B1(_05059_),
    .B2(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__or2_2 _19366_ (.A(_05058_),
    .B(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__a21bo_2 _19367_ (.A1(_05058_),
    .A2(_05065_),
    .B1_N(_05066_),
    .X(_05067_));
 sky130_fd_sc_hd__o21ba_2 _19368_ (.A1(_05016_),
    .A2(_05018_),
    .B1_N(_05012_),
    .X(_05068_));
 sky130_fd_sc_hd__buf_1 _19369_ (.A(_04706_),
    .X(_05069_));
 sky130_fd_sc_hd__buf_1 _19370_ (.A(_05014_),
    .X(_05070_));
 sky130_fd_sc_hd__buf_1 _19371_ (.A(_05020_),
    .X(_05071_));
 sky130_fd_sc_hd__buf_1 _19372_ (.A(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__o22a_2 _19373_ (.A1(_05069_),
    .A2(_05070_),
    .B1(_04693_),
    .B2(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__and4_2 _19374_ (.A(_11635_),
    .B(_11929_),
    .C(_11641_),
    .D(_11927_),
    .X(_05074_));
 sky130_fd_sc_hd__nor2_2 _19375_ (.A(_05073_),
    .B(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__buf_1 _19376_ (.A(_05013_),
    .X(_05076_));
 sky130_fd_sc_hd__buf_1 _19377_ (.A(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__nor2_2 _19378_ (.A(_04730_),
    .B(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__a2bb2o_2 _19379_ (.A1_N(_05075_),
    .A2_N(_05078_),
    .B1(_05075_),
    .B2(_05078_),
    .X(_05079_));
 sky130_vsdinv _19380_ (.A(\pcpi_mul.rs1[12] ),
    .Y(_05080_));
 sky130_fd_sc_hd__buf_1 _19381_ (.A(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__or2_2 _19382_ (.A(_04536_),
    .B(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__buf_1 _19383_ (.A(_04774_),
    .X(_05083_));
 sky130_fd_sc_hd__buf_1 _19384_ (.A(_04844_),
    .X(_05084_));
 sky130_fd_sc_hd__buf_1 _19385_ (.A(_04740_),
    .X(_05085_));
 sky130_fd_sc_hd__buf_1 _19386_ (.A(_04958_),
    .X(_05086_));
 sky130_fd_sc_hd__o22a_2 _19387_ (.A1(_05083_),
    .A2(_05084_),
    .B1(_05085_),
    .B2(_05086_),
    .X(_05087_));
 sky130_fd_sc_hd__and4_2 _19388_ (.A(_11626_),
    .B(_11936_),
    .C(_11630_),
    .D(_11933_),
    .X(_05088_));
 sky130_fd_sc_hd__or2_2 _19389_ (.A(_05087_),
    .B(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__a2bb2o_2 _19390_ (.A1_N(_05082_),
    .A2_N(_05089_),
    .B1(_05082_),
    .B2(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__o21ba_2 _19391_ (.A1(_05021_),
    .A2(_05024_),
    .B1_N(_05022_),
    .X(_05091_));
 sky130_fd_sc_hd__a2bb2o_2 _19392_ (.A1_N(_05090_),
    .A2_N(_05091_),
    .B1(_05090_),
    .B2(_05091_),
    .X(_05092_));
 sky130_fd_sc_hd__a2bb2o_2 _19393_ (.A1_N(_05079_),
    .A2_N(_05092_),
    .B1(_05079_),
    .B2(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__o22a_2 _19394_ (.A1(_05025_),
    .A2(_05026_),
    .B1(_05019_),
    .B2(_05027_),
    .X(_05094_));
 sky130_fd_sc_hd__a2bb2o_2 _19395_ (.A1_N(_05093_),
    .A2_N(_05094_),
    .B1(_05093_),
    .B2(_05094_),
    .X(_05095_));
 sky130_fd_sc_hd__a2bb2o_2 _19396_ (.A1_N(_05068_),
    .A2_N(_05095_),
    .B1(_05068_),
    .B2(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__or2_2 _19397_ (.A(_04983_),
    .B(_05039_),
    .X(_05097_));
 sky130_fd_sc_hd__o21ba_2 _19398_ (.A1(_05033_),
    .A2(_05036_),
    .B1_N(_05035_),
    .X(_05098_));
 sky130_fd_sc_hd__o21ba_2 _19399_ (.A1(_05005_),
    .A2(_05009_),
    .B1_N(_05006_),
    .X(_05099_));
 sky130_fd_sc_hd__buf_1 _19400_ (.A(_04807_),
    .X(_05100_));
 sky130_fd_sc_hd__or2_2 _19401_ (.A(_04793_),
    .B(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__o22a_2 _19402_ (.A1(_04977_),
    .A2(_04745_),
    .B1(_04826_),
    .B2(_04770_),
    .X(_05102_));
 sky130_fd_sc_hd__and4_2 _19403_ (.A(_11618_),
    .B(_11944_),
    .C(_11622_),
    .D(_11941_),
    .X(_05103_));
 sky130_fd_sc_hd__or2_2 _19404_ (.A(_05102_),
    .B(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__a2bb2o_2 _19405_ (.A1_N(_05101_),
    .A2_N(_05104_),
    .B1(_05101_),
    .B2(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__a2bb2o_2 _19406_ (.A1_N(_05099_),
    .A2_N(_05105_),
    .B1(_05099_),
    .B2(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__a2bb2o_2 _19407_ (.A1_N(_05098_),
    .A2_N(_05106_),
    .B1(_05098_),
    .B2(_05106_),
    .X(_05107_));
 sky130_fd_sc_hd__o22a_2 _19408_ (.A1(_04954_),
    .A2(_05037_),
    .B1(_05032_),
    .B2(_05038_),
    .X(_05108_));
 sky130_fd_sc_hd__or2_2 _19409_ (.A(_05107_),
    .B(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__a21bo_2 _19410_ (.A1(_05107_),
    .A2(_05108_),
    .B1_N(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__a2bb2o_2 _19411_ (.A1_N(_05097_),
    .A2_N(_05110_),
    .B1(_05097_),
    .B2(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__a2bb2o_2 _19412_ (.A1_N(_05096_),
    .A2_N(_05111_),
    .B1(_05096_),
    .B2(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__o32a_2 _19413_ (.A1(_04911_),
    .A2(_04984_),
    .A3(_05039_),
    .B1(_05031_),
    .B2(_05041_),
    .X(_05113_));
 sky130_fd_sc_hd__or2_2 _19414_ (.A(_05112_),
    .B(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__a21bo_2 _19415_ (.A1(_05112_),
    .A2(_05113_),
    .B1_N(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__or2_2 _19416_ (.A(_05067_),
    .B(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__a21bo_2 _19417_ (.A1(_05067_),
    .A2(_05115_),
    .B1_N(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__a2bb2o_2 _19418_ (.A1_N(_05046_),
    .A2_N(_05117_),
    .B1(_05046_),
    .B2(_05117_),
    .X(_05118_));
 sky130_fd_sc_hd__o22a_2 _19419_ (.A1(_05028_),
    .A2(_05029_),
    .B1(_05011_),
    .B2(_05030_),
    .X(_05119_));
 sky130_fd_sc_hd__or2_2 _19420_ (.A(_05044_),
    .B(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__a21bo_2 _19421_ (.A1(_05044_),
    .A2(_05119_),
    .B1_N(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__a2bb2o_2 _19422_ (.A1_N(_05118_),
    .A2_N(_05121_),
    .B1(_05118_),
    .B2(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__o22a_2 _19423_ (.A1(_04990_),
    .A2(_05047_),
    .B1(_05004_),
    .B2(_05048_),
    .X(_05123_));
 sky130_fd_sc_hd__a2bb2o_2 _19424_ (.A1_N(_05122_),
    .A2_N(_05123_),
    .B1(_05122_),
    .B2(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__a2bb2o_2 _19425_ (.A1_N(_05003_),
    .A2_N(_05124_),
    .B1(_05003_),
    .B2(_05124_),
    .X(_05125_));
 sky130_fd_sc_hd__o22a_2 _19426_ (.A1(_05049_),
    .A2(_05050_),
    .B1(_04994_),
    .B2(_05051_),
    .X(_05126_));
 sky130_fd_sc_hd__a2bb2o_2 _19427_ (.A1_N(_05125_),
    .A2_N(_05126_),
    .B1(_05125_),
    .B2(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__o22a_2 _19428_ (.A1(_04998_),
    .A2(_05052_),
    .B1(_05053_),
    .B2(_05054_),
    .X(_05128_));
 sky130_fd_sc_hd__a2bb2oi_2 _19429_ (.A1_N(_05127_),
    .A2_N(_05128_),
    .B1(_05127_),
    .B2(_05128_),
    .Y(_02631_));
 sky130_fd_sc_hd__o22a_2 _19430_ (.A1(_05125_),
    .A2(_05126_),
    .B1(_05127_),
    .B2(_05128_),
    .X(_05129_));
 sky130_vsdinv _19431_ (.A(\pcpi_mul.rs2[13] ),
    .Y(_05130_));
 sky130_fd_sc_hd__buf_1 _19432_ (.A(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__buf_1 _19433_ (.A(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__buf_1 _19434_ (.A(_05055_),
    .X(_05133_));
 sky130_fd_sc_hd__o22a_2 _19435_ (.A1(_05132_),
    .A2(_04707_),
    .B1(_05133_),
    .B2(_04689_),
    .X(_05134_));
 sky130_fd_sc_hd__or4_2 _19436_ (.A(_05132_),
    .B(_04707_),
    .C(_05056_),
    .D(_04703_),
    .X(_05135_));
 sky130_fd_sc_hd__or2b_2 _19437_ (.A(_05134_),
    .B_N(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__buf_1 _19438_ (.A(_04742_),
    .X(_05137_));
 sky130_fd_sc_hd__or2_2 _19439_ (.A(_04953_),
    .B(_05137_),
    .X(_05138_));
 sky130_fd_sc_hd__buf_1 _19440_ (.A(_05007_),
    .X(_05139_));
 sky130_fd_sc_hd__buf_1 _19441_ (.A(_04949_),
    .X(_05140_));
 sky130_fd_sc_hd__buf_1 _19442_ (.A(_04782_),
    .X(_05141_));
 sky130_fd_sc_hd__o22a_2 _19443_ (.A1(_05139_),
    .A2(_04701_),
    .B1(_05140_),
    .B2(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__buf_1 _19444_ (.A(\pcpi_mul.rs2[11] ),
    .X(_05143_));
 sky130_fd_sc_hd__buf_1 _19445_ (.A(_11951_),
    .X(_05144_));
 sky130_fd_sc_hd__buf_1 _19446_ (.A(_11947_),
    .X(_05145_));
 sky130_fd_sc_hd__and4_2 _19447_ (.A(_05143_),
    .B(_05144_),
    .C(_11615_),
    .D(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__or2_2 _19448_ (.A(_05142_),
    .B(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__a2bb2o_2 _19449_ (.A1_N(_05138_),
    .A2_N(_05147_),
    .B1(_05138_),
    .B2(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__or2_2 _19450_ (.A(_05136_),
    .B(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__a21bo_2 _19451_ (.A1(_05136_),
    .A2(_05148_),
    .B1_N(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__o22a_2 _19452_ (.A1(_05097_),
    .A2(_05110_),
    .B1(_05096_),
    .B2(_05111_),
    .X(_05151_));
 sky130_fd_sc_hd__a21oi_2 _19453_ (.A1(_05075_),
    .A2(_05078_),
    .B1(_05074_),
    .Y(_05152_));
 sky130_fd_sc_hd__buf_1 _19454_ (.A(_04706_),
    .X(_05153_));
 sky130_fd_sc_hd__buf_1 _19455_ (.A(_05071_),
    .X(_05154_));
 sky130_fd_sc_hd__buf_1 _19456_ (.A(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__buf_1 _19457_ (.A(_04693_),
    .X(_05156_));
 sky130_fd_sc_hd__buf_1 _19458_ (.A(_05080_),
    .X(_05157_));
 sky130_fd_sc_hd__buf_1 _19459_ (.A(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__o22a_2 _19460_ (.A1(_05153_),
    .A2(_05155_),
    .B1(_05156_),
    .B2(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__and4_2 _19461_ (.A(_11637_),
    .B(_11927_),
    .C(_11643_),
    .D(_11925_),
    .X(_05160_));
 sky130_fd_sc_hd__nor2_2 _19462_ (.A(_05159_),
    .B(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__buf_1 _19463_ (.A(_04730_),
    .X(_05162_));
 sky130_fd_sc_hd__buf_1 _19464_ (.A(_04963_),
    .X(_05163_));
 sky130_fd_sc_hd__buf_1 _19465_ (.A(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__nor2_2 _19466_ (.A(_05162_),
    .B(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__a2bb2o_2 _19467_ (.A1_N(_05161_),
    .A2_N(_05165_),
    .B1(_05161_),
    .B2(_05165_),
    .X(_05166_));
 sky130_vsdinv _19468_ (.A(\pcpi_mul.rs1[13] ),
    .Y(_05167_));
 sky130_fd_sc_hd__buf_1 _19469_ (.A(_05167_),
    .X(_05168_));
 sky130_fd_sc_hd__buf_1 _19470_ (.A(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__or2_2 _19471_ (.A(_04719_),
    .B(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__buf_1 _19472_ (.A(_05083_),
    .X(_05171_));
 sky130_fd_sc_hd__buf_1 _19473_ (.A(_04958_),
    .X(_05172_));
 sky130_fd_sc_hd__buf_1 _19474_ (.A(_05085_),
    .X(_05173_));
 sky130_fd_sc_hd__buf_1 _19475_ (.A(_05013_),
    .X(_05174_));
 sky130_fd_sc_hd__o22a_2 _19476_ (.A1(_05171_),
    .A2(_05172_),
    .B1(_05173_),
    .B2(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__buf_1 _19477_ (.A(_11933_),
    .X(_05176_));
 sky130_fd_sc_hd__buf_1 _19478_ (.A(\pcpi_mul.rs1[9] ),
    .X(_05177_));
 sky130_fd_sc_hd__and4_2 _19479_ (.A(_11627_),
    .B(_05176_),
    .C(_11631_),
    .D(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__or2_2 _19480_ (.A(_05175_),
    .B(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__a2bb2o_2 _19481_ (.A1_N(_05170_),
    .A2_N(_05179_),
    .B1(_05170_),
    .B2(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__o21ba_2 _19482_ (.A1(_05082_),
    .A2(_05089_),
    .B1_N(_05088_),
    .X(_05181_));
 sky130_fd_sc_hd__a2bb2o_2 _19483_ (.A1_N(_05180_),
    .A2_N(_05181_),
    .B1(_05180_),
    .B2(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__a2bb2o_2 _19484_ (.A1_N(_05166_),
    .A2_N(_05182_),
    .B1(_05166_),
    .B2(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__o22a_2 _19485_ (.A1(_05090_),
    .A2(_05091_),
    .B1(_05079_),
    .B2(_05092_),
    .X(_05184_));
 sky130_fd_sc_hd__a2bb2o_2 _19486_ (.A1_N(_05183_),
    .A2_N(_05184_),
    .B1(_05183_),
    .B2(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__a2bb2o_2 _19487_ (.A1_N(_05152_),
    .A2_N(_05185_),
    .B1(_05152_),
    .B2(_05185_),
    .X(_05186_));
 sky130_fd_sc_hd__o22a_2 _19488_ (.A1(_05099_),
    .A2(_05105_),
    .B1(_05098_),
    .B2(_05106_),
    .X(_05187_));
 sky130_fd_sc_hd__o21ba_2 _19489_ (.A1(_05101_),
    .A2(_05104_),
    .B1_N(_05103_),
    .X(_05188_));
 sky130_fd_sc_hd__o21ba_2 _19490_ (.A1(_05059_),
    .A2(_05064_),
    .B1_N(_05063_),
    .X(_05189_));
 sky130_fd_sc_hd__buf_1 _19491_ (.A(_04844_),
    .X(_05190_));
 sky130_fd_sc_hd__buf_1 _19492_ (.A(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__or2_2 _19493_ (.A(_04794_),
    .B(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__buf_1 _19494_ (.A(_04977_),
    .X(_05193_));
 sky130_fd_sc_hd__buf_1 _19495_ (.A(_04876_),
    .X(_05194_));
 sky130_fd_sc_hd__buf_1 _19496_ (.A(_05100_),
    .X(_05195_));
 sky130_fd_sc_hd__o22a_2 _19497_ (.A1(_05193_),
    .A2(_05194_),
    .B1(_04827_),
    .B2(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__buf_1 _19498_ (.A(_11941_),
    .X(_05197_));
 sky130_fd_sc_hd__buf_1 _19499_ (.A(_11938_),
    .X(_05198_));
 sky130_fd_sc_hd__and4_2 _19500_ (.A(_11619_),
    .B(_05197_),
    .C(_11623_),
    .D(_05198_),
    .X(_05199_));
 sky130_fd_sc_hd__or2_2 _19501_ (.A(_05196_),
    .B(_05199_),
    .X(_05200_));
 sky130_fd_sc_hd__a2bb2o_2 _19502_ (.A1_N(_05192_),
    .A2_N(_05200_),
    .B1(_05192_),
    .B2(_05200_),
    .X(_05201_));
 sky130_fd_sc_hd__a2bb2o_2 _19503_ (.A1_N(_05189_),
    .A2_N(_05201_),
    .B1(_05189_),
    .B2(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__a2bb2o_2 _19504_ (.A1_N(_05188_),
    .A2_N(_05202_),
    .B1(_05188_),
    .B2(_05202_),
    .X(_05203_));
 sky130_fd_sc_hd__a2bb2o_2 _19505_ (.A1_N(_05066_),
    .A2_N(_05203_),
    .B1(_05066_),
    .B2(_05203_),
    .X(_05204_));
 sky130_fd_sc_hd__a2bb2o_2 _19506_ (.A1_N(_05187_),
    .A2_N(_05204_),
    .B1(_05187_),
    .B2(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__a2bb2o_2 _19507_ (.A1_N(_05109_),
    .A2_N(_05205_),
    .B1(_05109_),
    .B2(_05205_),
    .X(_05206_));
 sky130_fd_sc_hd__a2bb2o_2 _19508_ (.A1_N(_05186_),
    .A2_N(_05206_),
    .B1(_05186_),
    .B2(_05206_),
    .X(_05207_));
 sky130_fd_sc_hd__or2_2 _19509_ (.A(_05151_),
    .B(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__a21bo_2 _19510_ (.A1(_05151_),
    .A2(_05207_),
    .B1_N(_05208_),
    .X(_05209_));
 sky130_fd_sc_hd__or2_2 _19511_ (.A(_05150_),
    .B(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__a21bo_2 _19512_ (.A1(_05150_),
    .A2(_05209_),
    .B1_N(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__a2bb2o_2 _19513_ (.A1_N(_05116_),
    .A2_N(_05211_),
    .B1(_05116_),
    .B2(_05211_),
    .X(_05212_));
 sky130_fd_sc_hd__o22a_2 _19514_ (.A1(_05093_),
    .A2(_05094_),
    .B1(_05068_),
    .B2(_05095_),
    .X(_05213_));
 sky130_fd_sc_hd__or2_2 _19515_ (.A(_05114_),
    .B(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__a21bo_2 _19516_ (.A1(_05114_),
    .A2(_05213_),
    .B1_N(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__a2bb2o_2 _19517_ (.A1_N(_05212_),
    .A2_N(_05215_),
    .B1(_05212_),
    .B2(_05215_),
    .X(_05216_));
 sky130_fd_sc_hd__o22a_2 _19518_ (.A1(_05046_),
    .A2(_05117_),
    .B1(_05118_),
    .B2(_05121_),
    .X(_05217_));
 sky130_fd_sc_hd__a2bb2o_2 _19519_ (.A1_N(_05216_),
    .A2_N(_05217_),
    .B1(_05216_),
    .B2(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__a2bb2o_2 _19520_ (.A1_N(_05120_),
    .A2_N(_05218_),
    .B1(_05120_),
    .B2(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__o22a_2 _19521_ (.A1(_05122_),
    .A2(_05123_),
    .B1(_05003_),
    .B2(_05124_),
    .X(_05220_));
 sky130_fd_sc_hd__a2bb2o_2 _19522_ (.A1_N(_05219_),
    .A2_N(_05220_),
    .B1(_05219_),
    .B2(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__a2bb2oi_2 _19523_ (.A1_N(_05129_),
    .A2_N(_05221_),
    .B1(_05129_),
    .B2(_05221_),
    .Y(_02632_));
 sky130_fd_sc_hd__o22a_2 _19524_ (.A1(_05183_),
    .A2(_05184_),
    .B1(_05152_),
    .B2(_05185_),
    .X(_05222_));
 sky130_fd_sc_hd__or2_2 _19525_ (.A(_05208_),
    .B(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__a21bo_2 _19526_ (.A1(_05208_),
    .A2(_05222_),
    .B1_N(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__buf_1 _19527_ (.A(_04876_),
    .X(_05225_));
 sky130_fd_sc_hd__or2_2 _19528_ (.A(_04953_),
    .B(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__buf_1 _19529_ (.A(_04745_),
    .X(_05227_));
 sky130_fd_sc_hd__o22a_2 _19530_ (.A1(_05139_),
    .A2(_04722_),
    .B1(_05140_),
    .B2(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__and4_2 _19531_ (.A(_05143_),
    .B(_05145_),
    .C(_11615_),
    .D(_11945_),
    .X(_05229_));
 sky130_fd_sc_hd__or2_2 _19532_ (.A(_05228_),
    .B(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__a2bb2o_2 _19533_ (.A1_N(_05226_),
    .A2_N(_05230_),
    .B1(_05226_),
    .B2(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__buf_1 _19534_ (.A(_05055_),
    .X(_05232_));
 sky130_fd_sc_hd__or2_2 _19535_ (.A(_05232_),
    .B(_04702_),
    .X(_05233_));
 sky130_vsdinv _19536_ (.A(\pcpi_mul.rs2[14] ),
    .Y(_05234_));
 sky130_fd_sc_hd__buf_1 _19537_ (.A(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__o22a_2 _19538_ (.A1(_05130_),
    .A2(_04709_),
    .B1(_05235_),
    .B2(_04710_),
    .X(_05236_));
 sky130_fd_sc_hd__buf_1 _19539_ (.A(\pcpi_mul.rs2[13] ),
    .X(_05237_));
 sky130_fd_sc_hd__buf_1 _19540_ (.A(_11953_),
    .X(_05238_));
 sky130_fd_sc_hd__and4_2 _19541_ (.A(_05237_),
    .B(_05238_),
    .C(\pcpi_mul.rs2[14] ),
    .D(_11957_),
    .X(_05239_));
 sky130_fd_sc_hd__or2_2 _19542_ (.A(_05236_),
    .B(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__a2bb2o_2 _19543_ (.A1_N(_05233_),
    .A2_N(_05240_),
    .B1(_05233_),
    .B2(_05240_),
    .X(_05241_));
 sky130_fd_sc_hd__a2bb2o_2 _19544_ (.A1_N(_05135_),
    .A2_N(_05241_),
    .B1(_05135_),
    .B2(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__a2bb2o_2 _19545_ (.A1_N(_05231_),
    .A2_N(_05242_),
    .B1(_05231_),
    .B2(_05242_),
    .X(_05243_));
 sky130_fd_sc_hd__o22a_2 _19546_ (.A1(_05109_),
    .A2(_05205_),
    .B1(_05186_),
    .B2(_05206_),
    .X(_05244_));
 sky130_fd_sc_hd__a21oi_2 _19547_ (.A1(_05161_),
    .A2(_05165_),
    .B1(_05160_),
    .Y(_05245_));
 sky130_fd_sc_hd__buf_1 _19548_ (.A(_05167_),
    .X(_05246_));
 sky130_fd_sc_hd__buf_1 _19549_ (.A(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__o22a_2 _19550_ (.A1(_05069_),
    .A2(_05158_),
    .B1(_04694_),
    .B2(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__and4_2 _19551_ (.A(_11636_),
    .B(_11925_),
    .C(_11642_),
    .D(_11923_),
    .X(_05249_));
 sky130_fd_sc_hd__nor2_2 _19552_ (.A(_05248_),
    .B(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__buf_1 _19553_ (.A(_04730_),
    .X(_05251_));
 sky130_fd_sc_hd__nor2_2 _19554_ (.A(_05251_),
    .B(_05155_),
    .Y(_05252_));
 sky130_fd_sc_hd__a2bb2o_2 _19555_ (.A1_N(_05250_),
    .A2_N(_05252_),
    .B1(_05250_),
    .B2(_05252_),
    .X(_05253_));
 sky130_vsdinv _19556_ (.A(\pcpi_mul.rs1[14] ),
    .Y(_05254_));
 sky130_fd_sc_hd__buf_1 _19557_ (.A(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__buf_1 _19558_ (.A(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__or2_2 _19559_ (.A(_04719_),
    .B(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__buf_1 _19560_ (.A(_05014_),
    .X(_05258_));
 sky130_fd_sc_hd__o22a_2 _19561_ (.A1(_05083_),
    .A2(_05174_),
    .B1(_05085_),
    .B2(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__buf_1 _19562_ (.A(\pcpi_mul.rs1[10] ),
    .X(_05260_));
 sky130_fd_sc_hd__and4_2 _19563_ (.A(_11627_),
    .B(_05177_),
    .C(_11631_),
    .D(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__or2_2 _19564_ (.A(_05259_),
    .B(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__a2bb2o_2 _19565_ (.A1_N(_05257_),
    .A2_N(_05262_),
    .B1(_05257_),
    .B2(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__o21ba_2 _19566_ (.A1(_05170_),
    .A2(_05179_),
    .B1_N(_05178_),
    .X(_05264_));
 sky130_fd_sc_hd__a2bb2o_2 _19567_ (.A1_N(_05263_),
    .A2_N(_05264_),
    .B1(_05263_),
    .B2(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__a2bb2o_2 _19568_ (.A1_N(_05253_),
    .A2_N(_05265_),
    .B1(_05253_),
    .B2(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__o22a_2 _19569_ (.A1(_05180_),
    .A2(_05181_),
    .B1(_05166_),
    .B2(_05182_),
    .X(_05267_));
 sky130_fd_sc_hd__a2bb2o_2 _19570_ (.A1_N(_05266_),
    .A2_N(_05267_),
    .B1(_05266_),
    .B2(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__a2bb2o_2 _19571_ (.A1_N(_05245_),
    .A2_N(_05268_),
    .B1(_05245_),
    .B2(_05268_),
    .X(_05269_));
 sky130_fd_sc_hd__o22a_2 _19572_ (.A1(_05189_),
    .A2(_05201_),
    .B1(_05188_),
    .B2(_05202_),
    .X(_05270_));
 sky130_fd_sc_hd__o21ba_2 _19573_ (.A1(_05192_),
    .A2(_05200_),
    .B1_N(_05199_),
    .X(_05271_));
 sky130_fd_sc_hd__o21ba_2 _19574_ (.A1(_05138_),
    .A2(_05147_),
    .B1_N(_05146_),
    .X(_05272_));
 sky130_fd_sc_hd__buf_1 _19575_ (.A(_04958_),
    .X(_05273_));
 sky130_fd_sc_hd__or2_2 _19576_ (.A(_04829_),
    .B(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__buf_1 _19577_ (.A(_04977_),
    .X(_05275_));
 sky130_fd_sc_hd__buf_1 _19578_ (.A(_04826_),
    .X(_05276_));
 sky130_fd_sc_hd__o22a_2 _19579_ (.A1(_05275_),
    .A2(_05100_),
    .B1(_05276_),
    .B2(_05084_),
    .X(_05277_));
 sky130_fd_sc_hd__buf_1 _19580_ (.A(_11618_),
    .X(_05278_));
 sky130_fd_sc_hd__buf_1 _19581_ (.A(_11622_),
    .X(_05279_));
 sky130_fd_sc_hd__buf_1 _19582_ (.A(_11936_),
    .X(_05280_));
 sky130_fd_sc_hd__and4_2 _19583_ (.A(_05278_),
    .B(_11939_),
    .C(_05279_),
    .D(_05280_),
    .X(_05281_));
 sky130_fd_sc_hd__or2_2 _19584_ (.A(_05277_),
    .B(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__a2bb2o_2 _19585_ (.A1_N(_05274_),
    .A2_N(_05282_),
    .B1(_05274_),
    .B2(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__a2bb2o_2 _19586_ (.A1_N(_05272_),
    .A2_N(_05283_),
    .B1(_05272_),
    .B2(_05283_),
    .X(_05284_));
 sky130_fd_sc_hd__a2bb2o_2 _19587_ (.A1_N(_05271_),
    .A2_N(_05284_),
    .B1(_05271_),
    .B2(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__a2bb2o_2 _19588_ (.A1_N(_05149_),
    .A2_N(_05285_),
    .B1(_05149_),
    .B2(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__a2bb2o_2 _19589_ (.A1_N(_05270_),
    .A2_N(_05286_),
    .B1(_05270_),
    .B2(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__o22a_2 _19590_ (.A1(_05066_),
    .A2(_05203_),
    .B1(_05187_),
    .B2(_05204_),
    .X(_05288_));
 sky130_fd_sc_hd__a2bb2o_2 _19591_ (.A1_N(_05287_),
    .A2_N(_05288_),
    .B1(_05287_),
    .B2(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__a2bb2o_2 _19592_ (.A1_N(_05269_),
    .A2_N(_05289_),
    .B1(_05269_),
    .B2(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__or2_2 _19593_ (.A(_05244_),
    .B(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__a21bo_2 _19594_ (.A1(_05244_),
    .A2(_05290_),
    .B1_N(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__or2_2 _19595_ (.A(_05243_),
    .B(_05292_),
    .X(_05293_));
 sky130_fd_sc_hd__a21bo_2 _19596_ (.A1(_05243_),
    .A2(_05292_),
    .B1_N(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__a2bb2o_2 _19597_ (.A1_N(_05210_),
    .A2_N(_05294_),
    .B1(_05210_),
    .B2(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__a2bb2o_2 _19598_ (.A1_N(_05224_),
    .A2_N(_05295_),
    .B1(_05224_),
    .B2(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__o22a_2 _19599_ (.A1(_05116_),
    .A2(_05211_),
    .B1(_05212_),
    .B2(_05215_),
    .X(_05297_));
 sky130_fd_sc_hd__a2bb2o_2 _19600_ (.A1_N(_05296_),
    .A2_N(_05297_),
    .B1(_05296_),
    .B2(_05297_),
    .X(_05298_));
 sky130_fd_sc_hd__a2bb2o_2 _19601_ (.A1_N(_05214_),
    .A2_N(_05298_),
    .B1(_05214_),
    .B2(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__o22a_2 _19602_ (.A1(_05216_),
    .A2(_05217_),
    .B1(_05120_),
    .B2(_05218_),
    .X(_05300_));
 sky130_fd_sc_hd__a2bb2o_2 _19603_ (.A1_N(_05299_),
    .A2_N(_05300_),
    .B1(_05299_),
    .B2(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__o22a_2 _19604_ (.A1(_05219_),
    .A2(_05220_),
    .B1(_05129_),
    .B2(_05221_),
    .X(_05302_));
 sky130_fd_sc_hd__a2bb2oi_2 _19605_ (.A1_N(_05301_),
    .A2_N(_05302_),
    .B1(_05301_),
    .B2(_05302_),
    .Y(_02633_));
 sky130_fd_sc_hd__o22a_2 _19606_ (.A1(_05299_),
    .A2(_05300_),
    .B1(_05301_),
    .B2(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__o22a_2 _19607_ (.A1(_05266_),
    .A2(_05267_),
    .B1(_05245_),
    .B2(_05268_),
    .X(_05304_));
 sky130_fd_sc_hd__or2_2 _19608_ (.A(_05291_),
    .B(_05304_),
    .X(_05305_));
 sky130_fd_sc_hd__a21bo_2 _19609_ (.A1(_05291_),
    .A2(_05304_),
    .B1_N(_05305_),
    .X(_05306_));
 sky130_vsdinv _19610_ (.A(\pcpi_mul.rs2[15] ),
    .Y(_05307_));
 sky130_fd_sc_hd__buf_1 _19611_ (.A(_05307_),
    .X(_05308_));
 sky130_fd_sc_hd__buf_1 _19612_ (.A(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__buf_1 _19613_ (.A(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__or2_2 _19614_ (.A(_05310_),
    .B(_04546_),
    .X(_05311_));
 sky130_fd_sc_hd__buf_1 _19615_ (.A(_05100_),
    .X(_05312_));
 sky130_fd_sc_hd__or2_2 _19616_ (.A(_04953_),
    .B(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__buf_1 _19617_ (.A(_04770_),
    .X(_05314_));
 sky130_fd_sc_hd__o22a_2 _19618_ (.A1(_05139_),
    .A2(_04975_),
    .B1(_05140_),
    .B2(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__buf_1 _19619_ (.A(_11944_),
    .X(_05316_));
 sky130_fd_sc_hd__and4_2 _19620_ (.A(_05143_),
    .B(_05316_),
    .C(_11615_),
    .D(_11942_),
    .X(_05317_));
 sky130_fd_sc_hd__or2_2 _19621_ (.A(_05315_),
    .B(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__a2bb2o_2 _19622_ (.A1_N(_05313_),
    .A2_N(_05318_),
    .B1(_05313_),
    .B2(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__or2_2 _19623_ (.A(_05232_),
    .B(_04723_),
    .X(_05320_));
 sky130_fd_sc_hd__buf_1 _19624_ (.A(_05130_),
    .X(_05321_));
 sky130_fd_sc_hd__o22a_2 _19625_ (.A1(_05235_),
    .A2(_04709_),
    .B1(_05321_),
    .B2(_04779_),
    .X(_05322_));
 sky130_fd_sc_hd__buf_1 _19626_ (.A(\pcpi_mul.rs2[14] ),
    .X(_05323_));
 sky130_fd_sc_hd__and4_2 _19627_ (.A(_05323_),
    .B(_05238_),
    .C(_05237_),
    .D(_05144_),
    .X(_05324_));
 sky130_fd_sc_hd__or2_2 _19628_ (.A(_05322_),
    .B(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__a2bb2o_2 _19629_ (.A1_N(_05320_),
    .A2_N(_05325_),
    .B1(_05320_),
    .B2(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__o21ba_2 _19630_ (.A1(_05233_),
    .A2(_05240_),
    .B1_N(_05239_),
    .X(_05327_));
 sky130_fd_sc_hd__a2bb2o_2 _19631_ (.A1_N(_05326_),
    .A2_N(_05327_),
    .B1(_05326_),
    .B2(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__a2bb2o_2 _19632_ (.A1_N(_05319_),
    .A2_N(_05328_),
    .B1(_05319_),
    .B2(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__nor2_2 _19633_ (.A(_05311_),
    .B(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__a21oi_2 _19634_ (.A1(_05311_),
    .A2(_05329_),
    .B1(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__o22a_2 _19635_ (.A1(_05287_),
    .A2(_05288_),
    .B1(_05269_),
    .B2(_05289_),
    .X(_05332_));
 sky130_fd_sc_hd__a21oi_2 _19636_ (.A1(_05250_),
    .A2(_05252_),
    .B1(_05249_),
    .Y(_05333_));
 sky130_fd_sc_hd__buf_1 _19637_ (.A(_05254_),
    .X(_05334_));
 sky130_fd_sc_hd__buf_1 _19638_ (.A(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__o22a_2 _19639_ (.A1(_05069_),
    .A2(_05247_),
    .B1(_04694_),
    .B2(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__and4_2 _19640_ (.A(_11636_),
    .B(_11923_),
    .C(_11642_),
    .D(_11920_),
    .X(_05337_));
 sky130_fd_sc_hd__nor2_2 _19641_ (.A(_05336_),
    .B(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__nor2_2 _19642_ (.A(_05251_),
    .B(_05158_),
    .Y(_05339_));
 sky130_fd_sc_hd__a2bb2o_2 _19643_ (.A1_N(_05338_),
    .A2_N(_05339_),
    .B1(_05338_),
    .B2(_05339_),
    .X(_05340_));
 sky130_vsdinv _19644_ (.A(\pcpi_mul.rs1[15] ),
    .Y(_05341_));
 sky130_fd_sc_hd__buf_1 _19645_ (.A(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__buf_1 _19646_ (.A(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__or2_2 _19647_ (.A(_04719_),
    .B(_05343_),
    .X(_05344_));
 sky130_fd_sc_hd__buf_1 _19648_ (.A(_05020_),
    .X(_05345_));
 sky130_fd_sc_hd__o22a_2 _19649_ (.A1(_05083_),
    .A2(_05163_),
    .B1(_05085_),
    .B2(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__and4_2 _19650_ (.A(_11627_),
    .B(_05260_),
    .C(_11631_),
    .D(_11926_),
    .X(_05347_));
 sky130_fd_sc_hd__or2_2 _19651_ (.A(_05346_),
    .B(_05347_),
    .X(_05348_));
 sky130_fd_sc_hd__a2bb2o_2 _19652_ (.A1_N(_05344_),
    .A2_N(_05348_),
    .B1(_05344_),
    .B2(_05348_),
    .X(_05349_));
 sky130_fd_sc_hd__o21ba_2 _19653_ (.A1(_05257_),
    .A2(_05262_),
    .B1_N(_05261_),
    .X(_05350_));
 sky130_fd_sc_hd__a2bb2o_2 _19654_ (.A1_N(_05349_),
    .A2_N(_05350_),
    .B1(_05349_),
    .B2(_05350_),
    .X(_05351_));
 sky130_fd_sc_hd__a2bb2o_2 _19655_ (.A1_N(_05340_),
    .A2_N(_05351_),
    .B1(_05340_),
    .B2(_05351_),
    .X(_05352_));
 sky130_fd_sc_hd__o22a_2 _19656_ (.A1(_05263_),
    .A2(_05264_),
    .B1(_05253_),
    .B2(_05265_),
    .X(_05353_));
 sky130_fd_sc_hd__a2bb2o_2 _19657_ (.A1_N(_05352_),
    .A2_N(_05353_),
    .B1(_05352_),
    .B2(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__a2bb2o_2 _19658_ (.A1_N(_05333_),
    .A2_N(_05354_),
    .B1(_05333_),
    .B2(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__o22a_2 _19659_ (.A1(_05272_),
    .A2(_05283_),
    .B1(_05271_),
    .B2(_05284_),
    .X(_05356_));
 sky130_fd_sc_hd__o22a_2 _19660_ (.A1(_05135_),
    .A2(_05241_),
    .B1(_05231_),
    .B2(_05242_),
    .X(_05357_));
 sky130_fd_sc_hd__o21ba_2 _19661_ (.A1(_05274_),
    .A2(_05282_),
    .B1_N(_05281_),
    .X(_05358_));
 sky130_fd_sc_hd__o21ba_2 _19662_ (.A1(_05226_),
    .A2(_05230_),
    .B1_N(_05229_),
    .X(_05359_));
 sky130_fd_sc_hd__or2_2 _19663_ (.A(_04829_),
    .B(_05174_),
    .X(_05360_));
 sky130_fd_sc_hd__o22a_2 _19664_ (.A1(_04977_),
    .A2(_05084_),
    .B1(_05276_),
    .B2(_05086_),
    .X(_05361_));
 sky130_fd_sc_hd__and4_2 _19665_ (.A(_05278_),
    .B(_11936_),
    .C(_05279_),
    .D(_11933_),
    .X(_05362_));
 sky130_fd_sc_hd__or2_2 _19666_ (.A(_05361_),
    .B(_05362_),
    .X(_05363_));
 sky130_fd_sc_hd__a2bb2o_2 _19667_ (.A1_N(_05360_),
    .A2_N(_05363_),
    .B1(_05360_),
    .B2(_05363_),
    .X(_05364_));
 sky130_fd_sc_hd__a2bb2o_2 _19668_ (.A1_N(_05359_),
    .A2_N(_05364_),
    .B1(_05359_),
    .B2(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__a2bb2o_2 _19669_ (.A1_N(_05358_),
    .A2_N(_05365_),
    .B1(_05358_),
    .B2(_05365_),
    .X(_05366_));
 sky130_fd_sc_hd__a2bb2o_2 _19670_ (.A1_N(_05357_),
    .A2_N(_05366_),
    .B1(_05357_),
    .B2(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__a2bb2o_2 _19671_ (.A1_N(_05356_),
    .A2_N(_05367_),
    .B1(_05356_),
    .B2(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__o22a_2 _19672_ (.A1(_05149_),
    .A2(_05285_),
    .B1(_05270_),
    .B2(_05286_),
    .X(_05369_));
 sky130_fd_sc_hd__a2bb2o_2 _19673_ (.A1_N(_05368_),
    .A2_N(_05369_),
    .B1(_05368_),
    .B2(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__a2bb2o_2 _19674_ (.A1_N(_05355_),
    .A2_N(_05370_),
    .B1(_05355_),
    .B2(_05370_),
    .X(_05371_));
 sky130_fd_sc_hd__or2_2 _19675_ (.A(_05332_),
    .B(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__a21boi_2 _19676_ (.A1(_05332_),
    .A2(_05371_),
    .B1_N(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__nand2_2 _19677_ (.A(_05331_),
    .B(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__o21ai_2 _19678_ (.A1(_05331_),
    .A2(_05373_),
    .B1(_05374_),
    .Y(_05375_));
 sky130_fd_sc_hd__a2bb2o_2 _19679_ (.A1_N(_05293_),
    .A2_N(_05375_),
    .B1(_05293_),
    .B2(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__a2bb2o_2 _19680_ (.A1_N(_05306_),
    .A2_N(_05376_),
    .B1(_05306_),
    .B2(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__o22a_2 _19681_ (.A1(_05210_),
    .A2(_05294_),
    .B1(_05224_),
    .B2(_05295_),
    .X(_05378_));
 sky130_fd_sc_hd__a2bb2o_2 _19682_ (.A1_N(_05377_),
    .A2_N(_05378_),
    .B1(_05377_),
    .B2(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__a2bb2o_2 _19683_ (.A1_N(_05223_),
    .A2_N(_05379_),
    .B1(_05223_),
    .B2(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__o22a_2 _19684_ (.A1(_05296_),
    .A2(_05297_),
    .B1(_05214_),
    .B2(_05298_),
    .X(_05381_));
 sky130_fd_sc_hd__a2bb2o_2 _19685_ (.A1_N(_05380_),
    .A2_N(_05381_),
    .B1(_05380_),
    .B2(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__a2bb2oi_2 _19686_ (.A1_N(_05303_),
    .A2_N(_05382_),
    .B1(_05303_),
    .B2(_05382_),
    .Y(_02634_));
 sky130_fd_sc_hd__o22a_2 _19687_ (.A1(_05380_),
    .A2(_05381_),
    .B1(_05303_),
    .B2(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__o22a_2 _19688_ (.A1(_05352_),
    .A2(_05353_),
    .B1(_05333_),
    .B2(_05354_),
    .X(_05384_));
 sky130_fd_sc_hd__or2_2 _19689_ (.A(_05372_),
    .B(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__a21bo_2 _19690_ (.A1(_05372_),
    .A2(_05384_),
    .B1_N(_05385_),
    .X(_05386_));
 sky130_vsdinv _19691_ (.A(\pcpi_mul.rs2[16] ),
    .Y(_05387_));
 sky130_fd_sc_hd__buf_1 _19692_ (.A(_05387_),
    .X(_05388_));
 sky130_fd_sc_hd__buf_1 _19693_ (.A(_05388_),
    .X(_05389_));
 sky130_fd_sc_hd__o22a_2 _19694_ (.A1(_05389_),
    .A2(_04545_),
    .B1(_05310_),
    .B2(_04690_),
    .X(_05390_));
 sky130_fd_sc_hd__buf_1 _19695_ (.A(_05387_),
    .X(_05391_));
 sky130_fd_sc_hd__buf_1 _19696_ (.A(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__buf_1 _19697_ (.A(_05307_),
    .X(_05393_));
 sky130_fd_sc_hd__or4_2 _19698_ (.A(_05392_),
    .B(_04707_),
    .C(_05393_),
    .D(_04703_),
    .X(_05394_));
 sky130_fd_sc_hd__or2b_2 _19699_ (.A(_05390_),
    .B_N(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__buf_1 _19700_ (.A(_05084_),
    .X(_05396_));
 sky130_fd_sc_hd__or2_2 _19701_ (.A(_04902_),
    .B(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__buf_1 _19702_ (.A(_04807_),
    .X(_05398_));
 sky130_fd_sc_hd__o22a_2 _19703_ (.A1(_05060_),
    .A2(_05314_),
    .B1(_04950_),
    .B2(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__and4_2 _19704_ (.A(_11613_),
    .B(_05197_),
    .C(_11616_),
    .D(_11939_),
    .X(_05400_));
 sky130_fd_sc_hd__or2_2 _19705_ (.A(_05399_),
    .B(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__a2bb2o_2 _19706_ (.A1_N(_05397_),
    .A2_N(_05401_),
    .B1(_05397_),
    .B2(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__buf_1 _19707_ (.A(_05227_),
    .X(_05403_));
 sky130_fd_sc_hd__or2_2 _19708_ (.A(_05056_),
    .B(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__buf_1 _19709_ (.A(_05234_),
    .X(_05405_));
 sky130_fd_sc_hd__buf_1 _19710_ (.A(_04782_),
    .X(_05406_));
 sky130_fd_sc_hd__o22a_2 _19711_ (.A1(_05405_),
    .A2(_05061_),
    .B1(_05321_),
    .B2(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__and4_2 _19712_ (.A(_05323_),
    .B(_11952_),
    .C(_05237_),
    .D(_05145_),
    .X(_05408_));
 sky130_fd_sc_hd__or2_2 _19713_ (.A(_05407_),
    .B(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__a2bb2o_2 _19714_ (.A1_N(_05404_),
    .A2_N(_05409_),
    .B1(_05404_),
    .B2(_05409_),
    .X(_05410_));
 sky130_fd_sc_hd__o21ba_2 _19715_ (.A1(_05320_),
    .A2(_05325_),
    .B1_N(_05324_),
    .X(_05411_));
 sky130_fd_sc_hd__a2bb2o_2 _19716_ (.A1_N(_05410_),
    .A2_N(_05411_),
    .B1(_05410_),
    .B2(_05411_),
    .X(_05412_));
 sky130_fd_sc_hd__a2bb2o_2 _19717_ (.A1_N(_05402_),
    .A2_N(_05412_),
    .B1(_05402_),
    .B2(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__nor2_2 _19718_ (.A(_05395_),
    .B(_05413_),
    .Y(_05414_));
 sky130_fd_sc_hd__a21oi_2 _19719_ (.A1(_05395_),
    .A2(_05413_),
    .B1(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hd__nand2_2 _19720_ (.A(_05330_),
    .B(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__o21ai_2 _19721_ (.A1(_05330_),
    .A2(_05415_),
    .B1(_05416_),
    .Y(_05417_));
 sky130_fd_sc_hd__o22a_2 _19722_ (.A1(_05368_),
    .A2(_05369_),
    .B1(_05355_),
    .B2(_05370_),
    .X(_05418_));
 sky130_fd_sc_hd__a21oi_2 _19723_ (.A1(_05338_),
    .A2(_05339_),
    .B1(_05337_),
    .Y(_05419_));
 sky130_fd_sc_hd__buf_1 _19724_ (.A(_05342_),
    .X(_05420_));
 sky130_fd_sc_hd__buf_1 _19725_ (.A(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__o22a_2 _19726_ (.A1(_05069_),
    .A2(_05335_),
    .B1(_04694_),
    .B2(_05421_),
    .X(_05422_));
 sky130_fd_sc_hd__and4_2 _19727_ (.A(_11636_),
    .B(_11920_),
    .C(_11642_),
    .D(_11917_),
    .X(_05423_));
 sky130_fd_sc_hd__nor2_2 _19728_ (.A(_05422_),
    .B(_05423_),
    .Y(_05424_));
 sky130_fd_sc_hd__nor2_2 _19729_ (.A(_05251_),
    .B(_05247_),
    .Y(_05425_));
 sky130_fd_sc_hd__a2bb2o_2 _19730_ (.A1_N(_05424_),
    .A2_N(_05425_),
    .B1(_05424_),
    .B2(_05425_),
    .X(_05426_));
 sky130_vsdinv _19731_ (.A(\pcpi_mul.rs1[16] ),
    .Y(_05427_));
 sky130_fd_sc_hd__buf_1 _19732_ (.A(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__buf_1 _19733_ (.A(_05428_),
    .X(_05429_));
 sky130_fd_sc_hd__or2_2 _19734_ (.A(_04719_),
    .B(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__buf_1 _19735_ (.A(_05080_),
    .X(_05431_));
 sky130_fd_sc_hd__o22a_2 _19736_ (.A1(_05083_),
    .A2(_05345_),
    .B1(_05085_),
    .B2(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__buf_1 _19737_ (.A(\pcpi_mul.rs1[11] ),
    .X(_05433_));
 sky130_fd_sc_hd__and4_2 _19738_ (.A(_11627_),
    .B(_05433_),
    .C(_11631_),
    .D(_11924_),
    .X(_05434_));
 sky130_fd_sc_hd__or2_2 _19739_ (.A(_05432_),
    .B(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__a2bb2o_2 _19740_ (.A1_N(_05430_),
    .A2_N(_05435_),
    .B1(_05430_),
    .B2(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__o21ba_2 _19741_ (.A1(_05344_),
    .A2(_05348_),
    .B1_N(_05347_),
    .X(_05437_));
 sky130_fd_sc_hd__a2bb2o_2 _19742_ (.A1_N(_05436_),
    .A2_N(_05437_),
    .B1(_05436_),
    .B2(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__a2bb2o_2 _19743_ (.A1_N(_05426_),
    .A2_N(_05438_),
    .B1(_05426_),
    .B2(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__o22a_2 _19744_ (.A1(_05349_),
    .A2(_05350_),
    .B1(_05340_),
    .B2(_05351_),
    .X(_05440_));
 sky130_fd_sc_hd__a2bb2o_2 _19745_ (.A1_N(_05439_),
    .A2_N(_05440_),
    .B1(_05439_),
    .B2(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__a2bb2o_2 _19746_ (.A1_N(_05419_),
    .A2_N(_05441_),
    .B1(_05419_),
    .B2(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__o22a_2 _19747_ (.A1(_05359_),
    .A2(_05364_),
    .B1(_05358_),
    .B2(_05365_),
    .X(_05443_));
 sky130_fd_sc_hd__o22a_2 _19748_ (.A1(_05326_),
    .A2(_05327_),
    .B1(_05319_),
    .B2(_05328_),
    .X(_05444_));
 sky130_fd_sc_hd__o21ba_2 _19749_ (.A1(_05360_),
    .A2(_05363_),
    .B1_N(_05362_),
    .X(_05445_));
 sky130_fd_sc_hd__o21ba_2 _19750_ (.A1(_05313_),
    .A2(_05318_),
    .B1_N(_05317_),
    .X(_05446_));
 sky130_fd_sc_hd__or2_2 _19751_ (.A(_04829_),
    .B(_05258_),
    .X(_05447_));
 sky130_fd_sc_hd__o22a_2 _19752_ (.A1(_05275_),
    .A2(_04958_),
    .B1(_05276_),
    .B2(_05013_),
    .X(_05448_));
 sky130_fd_sc_hd__and4_2 _19753_ (.A(_05278_),
    .B(_11933_),
    .C(_05279_),
    .D(_11930_),
    .X(_05449_));
 sky130_fd_sc_hd__or2_2 _19754_ (.A(_05448_),
    .B(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__a2bb2o_2 _19755_ (.A1_N(_05447_),
    .A2_N(_05450_),
    .B1(_05447_),
    .B2(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__a2bb2o_2 _19756_ (.A1_N(_05446_),
    .A2_N(_05451_),
    .B1(_05446_),
    .B2(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__a2bb2o_2 _19757_ (.A1_N(_05445_),
    .A2_N(_05452_),
    .B1(_05445_),
    .B2(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__a2bb2o_2 _19758_ (.A1_N(_05444_),
    .A2_N(_05453_),
    .B1(_05444_),
    .B2(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__a2bb2o_2 _19759_ (.A1_N(_05443_),
    .A2_N(_05454_),
    .B1(_05443_),
    .B2(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__o22a_2 _19760_ (.A1(_05357_),
    .A2(_05366_),
    .B1(_05356_),
    .B2(_05367_),
    .X(_05456_));
 sky130_fd_sc_hd__a2bb2o_2 _19761_ (.A1_N(_05455_),
    .A2_N(_05456_),
    .B1(_05455_),
    .B2(_05456_),
    .X(_05457_));
 sky130_fd_sc_hd__a2bb2o_2 _19762_ (.A1_N(_05442_),
    .A2_N(_05457_),
    .B1(_05442_),
    .B2(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__or2_2 _19763_ (.A(_05418_),
    .B(_05458_),
    .X(_05459_));
 sky130_fd_sc_hd__a21bo_2 _19764_ (.A1(_05418_),
    .A2(_05458_),
    .B1_N(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__or2_2 _19765_ (.A(_05417_),
    .B(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__a21bo_2 _19766_ (.A1(_05417_),
    .A2(_05460_),
    .B1_N(_05461_),
    .X(_05462_));
 sky130_fd_sc_hd__a2bb2o_2 _19767_ (.A1_N(_05374_),
    .A2_N(_05462_),
    .B1(_05374_),
    .B2(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__a2bb2o_2 _19768_ (.A1_N(_05386_),
    .A2_N(_05463_),
    .B1(_05386_),
    .B2(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__o22a_2 _19769_ (.A1(_05293_),
    .A2(_05375_),
    .B1(_05306_),
    .B2(_05376_),
    .X(_05465_));
 sky130_fd_sc_hd__a2bb2o_2 _19770_ (.A1_N(_05464_),
    .A2_N(_05465_),
    .B1(_05464_),
    .B2(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__a2bb2o_2 _19771_ (.A1_N(_05305_),
    .A2_N(_05466_),
    .B1(_05305_),
    .B2(_05466_),
    .X(_05467_));
 sky130_fd_sc_hd__o22a_2 _19772_ (.A1(_05377_),
    .A2(_05378_),
    .B1(_05223_),
    .B2(_05379_),
    .X(_05468_));
 sky130_fd_sc_hd__or2_2 _19773_ (.A(_05467_),
    .B(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__a21bo_2 _19774_ (.A1(_05467_),
    .A2(_05468_),
    .B1_N(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__a2bb2oi_2 _19775_ (.A1_N(_05383_),
    .A2_N(_05470_),
    .B1(_05383_),
    .B2(_05470_),
    .Y(_02635_));
 sky130_fd_sc_hd__o22a_2 _19776_ (.A1(_05439_),
    .A2(_05440_),
    .B1(_05419_),
    .B2(_05441_),
    .X(_05471_));
 sky130_fd_sc_hd__or2_2 _19777_ (.A(_05459_),
    .B(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__a21bo_2 _19778_ (.A1(_05459_),
    .A2(_05471_),
    .B1_N(_05472_),
    .X(_05473_));
 sky130_fd_sc_hd__or2_2 _19779_ (.A(_05307_),
    .B(_04701_),
    .X(_05474_));
 sky130_vsdinv _19780_ (.A(\pcpi_mul.rs2[17] ),
    .Y(_05475_));
 sky130_fd_sc_hd__o22a_2 _19781_ (.A1(_05387_),
    .A2(_04686_),
    .B1(_05475_),
    .B2(_04541_),
    .X(_05476_));
 sky130_fd_sc_hd__and4_2 _19782_ (.A(_11604_),
    .B(_11954_),
    .C(\pcpi_mul.rs2[17] ),
    .D(_11956_),
    .X(_05477_));
 sky130_fd_sc_hd__or2_2 _19783_ (.A(_05476_),
    .B(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__a2bb2o_2 _19784_ (.A1_N(_05474_),
    .A2_N(_05478_),
    .B1(_05474_),
    .B2(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__or2_2 _19785_ (.A(_05394_),
    .B(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__a21bo_2 _19786_ (.A1(_05394_),
    .A2(_05479_),
    .B1_N(_05480_),
    .X(_05481_));
 sky130_fd_sc_hd__or2_2 _19787_ (.A(_04953_),
    .B(_05017_),
    .X(_05482_));
 sky130_fd_sc_hd__o22a_2 _19788_ (.A1(_05139_),
    .A2(_05398_),
    .B1(_05140_),
    .B2(_05084_),
    .X(_05483_));
 sky130_fd_sc_hd__and4_2 _19789_ (.A(_05143_),
    .B(_11939_),
    .C(_11615_),
    .D(_05280_),
    .X(_05484_));
 sky130_fd_sc_hd__or2_2 _19790_ (.A(_05483_),
    .B(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__a2bb2o_2 _19791_ (.A1_N(_05482_),
    .A2_N(_05485_),
    .B1(_05482_),
    .B2(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__or2_2 _19792_ (.A(_05232_),
    .B(_05225_),
    .X(_05487_));
 sky130_fd_sc_hd__o22a_2 _19793_ (.A1(_05235_),
    .A2(_04722_),
    .B1(_05321_),
    .B2(_04975_),
    .X(_05488_));
 sky130_fd_sc_hd__and4_2 _19794_ (.A(_05323_),
    .B(_11948_),
    .C(_05237_),
    .D(_11945_),
    .X(_05489_));
 sky130_fd_sc_hd__or2_2 _19795_ (.A(_05488_),
    .B(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__a2bb2o_2 _19796_ (.A1_N(_05487_),
    .A2_N(_05490_),
    .B1(_05487_),
    .B2(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__o21ba_2 _19797_ (.A1(_05404_),
    .A2(_05409_),
    .B1_N(_05408_),
    .X(_05492_));
 sky130_fd_sc_hd__a2bb2o_2 _19798_ (.A1_N(_05491_),
    .A2_N(_05492_),
    .B1(_05491_),
    .B2(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__a2bb2o_2 _19799_ (.A1_N(_05486_),
    .A2_N(_05493_),
    .B1(_05486_),
    .B2(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__nor2_2 _19800_ (.A(_05481_),
    .B(_05494_),
    .Y(_05495_));
 sky130_fd_sc_hd__a21oi_2 _19801_ (.A1(_05481_),
    .A2(_05494_),
    .B1(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__nand2_2 _19802_ (.A(_05414_),
    .B(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__o21ai_2 _19803_ (.A1(_05414_),
    .A2(_05496_),
    .B1(_05497_),
    .Y(_05498_));
 sky130_fd_sc_hd__o22a_2 _19804_ (.A1(_05455_),
    .A2(_05456_),
    .B1(_05442_),
    .B2(_05457_),
    .X(_05499_));
 sky130_fd_sc_hd__a21oi_2 _19805_ (.A1(_05424_),
    .A2(_05425_),
    .B1(_05423_),
    .Y(_05500_));
 sky130_fd_sc_hd__buf_1 _19806_ (.A(_05427_),
    .X(_05501_));
 sky130_fd_sc_hd__buf_1 _19807_ (.A(_05501_),
    .X(_05502_));
 sky130_fd_sc_hd__o22a_2 _19808_ (.A1(_05153_),
    .A2(_05421_),
    .B1(_05156_),
    .B2(_05502_),
    .X(_05503_));
 sky130_fd_sc_hd__and4_2 _19809_ (.A(_11637_),
    .B(_11917_),
    .C(_11643_),
    .D(_11915_),
    .X(_05504_));
 sky130_fd_sc_hd__nor2_2 _19810_ (.A(_05503_),
    .B(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__nor2_2 _19811_ (.A(_05251_),
    .B(_05335_),
    .Y(_05506_));
 sky130_fd_sc_hd__a2bb2o_2 _19812_ (.A1_N(_05505_),
    .A2_N(_05506_),
    .B1(_05505_),
    .B2(_05506_),
    .X(_05507_));
 sky130_vsdinv _19813_ (.A(\pcpi_mul.rs1[17] ),
    .Y(_05508_));
 sky130_fd_sc_hd__buf_1 _19814_ (.A(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__buf_1 _19815_ (.A(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__or2_2 _19816_ (.A(_04537_),
    .B(_05510_),
    .X(_05511_));
 sky130_fd_sc_hd__o22a_2 _19817_ (.A1(_05171_),
    .A2(_05431_),
    .B1(_05173_),
    .B2(_05246_),
    .X(_05512_));
 sky130_fd_sc_hd__buf_1 _19818_ (.A(_11627_),
    .X(_05513_));
 sky130_fd_sc_hd__buf_1 _19819_ (.A(\pcpi_mul.rs1[12] ),
    .X(_05514_));
 sky130_fd_sc_hd__buf_1 _19820_ (.A(_11631_),
    .X(_05515_));
 sky130_fd_sc_hd__buf_1 _19821_ (.A(\pcpi_mul.rs1[13] ),
    .X(_05516_));
 sky130_fd_sc_hd__and4_2 _19822_ (.A(_05513_),
    .B(_05514_),
    .C(_05515_),
    .D(_05516_),
    .X(_05517_));
 sky130_fd_sc_hd__or2_2 _19823_ (.A(_05512_),
    .B(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__a2bb2o_2 _19824_ (.A1_N(_05511_),
    .A2_N(_05518_),
    .B1(_05511_),
    .B2(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__o21ba_2 _19825_ (.A1(_05430_),
    .A2(_05435_),
    .B1_N(_05434_),
    .X(_05520_));
 sky130_fd_sc_hd__a2bb2o_2 _19826_ (.A1_N(_05519_),
    .A2_N(_05520_),
    .B1(_05519_),
    .B2(_05520_),
    .X(_05521_));
 sky130_fd_sc_hd__a2bb2o_2 _19827_ (.A1_N(_05507_),
    .A2_N(_05521_),
    .B1(_05507_),
    .B2(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__o22a_2 _19828_ (.A1(_05436_),
    .A2(_05437_),
    .B1(_05426_),
    .B2(_05438_),
    .X(_05523_));
 sky130_fd_sc_hd__a2bb2o_2 _19829_ (.A1_N(_05522_),
    .A2_N(_05523_),
    .B1(_05522_),
    .B2(_05523_),
    .X(_05524_));
 sky130_fd_sc_hd__a2bb2o_2 _19830_ (.A1_N(_05500_),
    .A2_N(_05524_),
    .B1(_05500_),
    .B2(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__o22a_2 _19831_ (.A1(_05446_),
    .A2(_05451_),
    .B1(_05445_),
    .B2(_05452_),
    .X(_05526_));
 sky130_fd_sc_hd__o22a_2 _19832_ (.A1(_05410_),
    .A2(_05411_),
    .B1(_05402_),
    .B2(_05412_),
    .X(_05527_));
 sky130_fd_sc_hd__o21ba_2 _19833_ (.A1(_05447_),
    .A2(_05450_),
    .B1_N(_05449_),
    .X(_05528_));
 sky130_fd_sc_hd__o21ba_2 _19834_ (.A1(_05397_),
    .A2(_05401_),
    .B1_N(_05400_),
    .X(_05529_));
 sky130_fd_sc_hd__buf_1 _19835_ (.A(_05071_),
    .X(_05530_));
 sky130_fd_sc_hd__or2_2 _19836_ (.A(_04794_),
    .B(_05530_),
    .X(_05531_));
 sky130_fd_sc_hd__o22a_2 _19837_ (.A1(_05275_),
    .A2(_05076_),
    .B1(_04827_),
    .B2(_05163_),
    .X(_05532_));
 sky130_fd_sc_hd__and4_2 _19838_ (.A(_05278_),
    .B(_11930_),
    .C(_05279_),
    .D(_11928_),
    .X(_05533_));
 sky130_fd_sc_hd__or2_2 _19839_ (.A(_05532_),
    .B(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__a2bb2o_2 _19840_ (.A1_N(_05531_),
    .A2_N(_05534_),
    .B1(_05531_),
    .B2(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__a2bb2o_2 _19841_ (.A1_N(_05529_),
    .A2_N(_05535_),
    .B1(_05529_),
    .B2(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__a2bb2o_2 _19842_ (.A1_N(_05528_),
    .A2_N(_05536_),
    .B1(_05528_),
    .B2(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__a2bb2o_2 _19843_ (.A1_N(_05527_),
    .A2_N(_05537_),
    .B1(_05527_),
    .B2(_05537_),
    .X(_05538_));
 sky130_fd_sc_hd__a2bb2o_2 _19844_ (.A1_N(_05526_),
    .A2_N(_05538_),
    .B1(_05526_),
    .B2(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__o22a_2 _19845_ (.A1(_05444_),
    .A2(_05453_),
    .B1(_05443_),
    .B2(_05454_),
    .X(_05540_));
 sky130_fd_sc_hd__a2bb2o_2 _19846_ (.A1_N(_05539_),
    .A2_N(_05540_),
    .B1(_05539_),
    .B2(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__a2bb2o_2 _19847_ (.A1_N(_05525_),
    .A2_N(_05541_),
    .B1(_05525_),
    .B2(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__a2bb2o_2 _19848_ (.A1_N(_05416_),
    .A2_N(_05542_),
    .B1(_05416_),
    .B2(_05542_),
    .X(_05543_));
 sky130_fd_sc_hd__a2bb2o_2 _19849_ (.A1_N(_05499_),
    .A2_N(_05543_),
    .B1(_05499_),
    .B2(_05543_),
    .X(_05544_));
 sky130_fd_sc_hd__or2_2 _19850_ (.A(_05498_),
    .B(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__a21bo_2 _19851_ (.A1(_05498_),
    .A2(_05544_),
    .B1_N(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__a2bb2o_2 _19852_ (.A1_N(_05461_),
    .A2_N(_05546_),
    .B1(_05461_),
    .B2(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__a2bb2o_2 _19853_ (.A1_N(_05473_),
    .A2_N(_05547_),
    .B1(_05473_),
    .B2(_05547_),
    .X(_05548_));
 sky130_fd_sc_hd__o22a_2 _19854_ (.A1(_05374_),
    .A2(_05462_),
    .B1(_05386_),
    .B2(_05463_),
    .X(_05549_));
 sky130_fd_sc_hd__a2bb2o_2 _19855_ (.A1_N(_05548_),
    .A2_N(_05549_),
    .B1(_05548_),
    .B2(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__a2bb2o_2 _19856_ (.A1_N(_05385_),
    .A2_N(_05550_),
    .B1(_05385_),
    .B2(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__o22a_2 _19857_ (.A1(_05464_),
    .A2(_05465_),
    .B1(_05305_),
    .B2(_05466_),
    .X(_05552_));
 sky130_fd_sc_hd__or2_2 _19858_ (.A(_05551_),
    .B(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__a21bo_2 _19859_ (.A1(_05551_),
    .A2(_05552_),
    .B1_N(_05553_),
    .X(_05554_));
 sky130_fd_sc_hd__o21ai_2 _19860_ (.A1(_05383_),
    .A2(_05470_),
    .B1(_05469_),
    .Y(_05555_));
 sky130_fd_sc_hd__a2bb2o_2 _19861_ (.A1_N(_05554_),
    .A2_N(_05555_),
    .B1(_05554_),
    .B2(_05555_),
    .X(_02636_));
 sky130_fd_sc_hd__o22a_2 _19862_ (.A1(_05416_),
    .A2(_05542_),
    .B1(_05499_),
    .B2(_05543_),
    .X(_05556_));
 sky130_fd_sc_hd__o22a_2 _19863_ (.A1(_05522_),
    .A2(_05523_),
    .B1(_05500_),
    .B2(_05524_),
    .X(_05557_));
 sky130_fd_sc_hd__or2_2 _19864_ (.A(_05556_),
    .B(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__a21bo_2 _19865_ (.A1(_05556_),
    .A2(_05557_),
    .B1_N(_05558_),
    .X(_05559_));
 sky130_vsdinv _19866_ (.A(\pcpi_mul.rs2[18] ),
    .Y(_05560_));
 sky130_fd_sc_hd__buf_1 _19867_ (.A(_05560_),
    .X(_05561_));
 sky130_fd_sc_hd__buf_1 _19868_ (.A(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__buf_1 _19869_ (.A(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__or2_2 _19870_ (.A(_05563_),
    .B(_04546_),
    .X(_05564_));
 sky130_fd_sc_hd__or2_2 _19871_ (.A(_05307_),
    .B(_04722_),
    .X(_05565_));
 sky130_fd_sc_hd__o22a_2 _19872_ (.A1(_05475_),
    .A2(_04686_),
    .B1(_05387_),
    .B2(_04699_),
    .X(_05566_));
 sky130_fd_sc_hd__and4_2 _19873_ (.A(\pcpi_mul.rs2[17] ),
    .B(_11953_),
    .C(\pcpi_mul.rs2[16] ),
    .D(_11950_),
    .X(_05567_));
 sky130_fd_sc_hd__or2_2 _19874_ (.A(_05566_),
    .B(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__a2bb2o_2 _19875_ (.A1_N(_05565_),
    .A2_N(_05568_),
    .B1(_05565_),
    .B2(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__o21ba_2 _19876_ (.A1(_05474_),
    .A2(_05478_),
    .B1_N(_05477_),
    .X(_05570_));
 sky130_fd_sc_hd__or2_2 _19877_ (.A(_05569_),
    .B(_05570_),
    .X(_05571_));
 sky130_fd_sc_hd__a21bo_2 _19878_ (.A1(_05569_),
    .A2(_05570_),
    .B1_N(_05571_),
    .X(_05572_));
 sky130_fd_sc_hd__o2bb2ai_2 _19879_ (.A1_N(_05480_),
    .A2_N(_05572_),
    .B1(_05480_),
    .B2(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__or2_2 _19880_ (.A(_04902_),
    .B(_05077_),
    .X(_05574_));
 sky130_fd_sc_hd__buf_1 _19881_ (.A(_04844_),
    .X(_05575_));
 sky130_fd_sc_hd__o22a_2 _19882_ (.A1(_05060_),
    .A2(_05575_),
    .B1(_04950_),
    .B2(_05273_),
    .X(_05576_));
 sky130_fd_sc_hd__buf_1 _19883_ (.A(_11936_),
    .X(_05577_));
 sky130_fd_sc_hd__buf_1 _19884_ (.A(_11933_),
    .X(_05578_));
 sky130_fd_sc_hd__and4_2 _19885_ (.A(_11613_),
    .B(_05577_),
    .C(_11616_),
    .D(_05578_),
    .X(_05579_));
 sky130_fd_sc_hd__or2_2 _19886_ (.A(_05576_),
    .B(_05579_),
    .X(_05580_));
 sky130_fd_sc_hd__a2bb2o_2 _19887_ (.A1_N(_05574_),
    .A2_N(_05580_),
    .B1(_05574_),
    .B2(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__or2_2 _19888_ (.A(_05232_),
    .B(_05195_),
    .X(_05582_));
 sky130_fd_sc_hd__o22a_2 _19889_ (.A1(_05235_),
    .A2(_04975_),
    .B1(_05130_),
    .B2(_05314_),
    .X(_05583_));
 sky130_fd_sc_hd__and4_2 _19890_ (.A(_05323_),
    .B(_11945_),
    .C(\pcpi_mul.rs2[13] ),
    .D(_11942_),
    .X(_05584_));
 sky130_fd_sc_hd__or2_2 _19891_ (.A(_05583_),
    .B(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__a2bb2o_2 _19892_ (.A1_N(_05582_),
    .A2_N(_05585_),
    .B1(_05582_),
    .B2(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__o21ba_2 _19893_ (.A1(_05487_),
    .A2(_05490_),
    .B1_N(_05489_),
    .X(_05587_));
 sky130_fd_sc_hd__a2bb2o_2 _19894_ (.A1_N(_05586_),
    .A2_N(_05587_),
    .B1(_05586_),
    .B2(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__a2bb2o_2 _19895_ (.A1_N(_05581_),
    .A2_N(_05588_),
    .B1(_05581_),
    .B2(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__o2bb2a_2 _19896_ (.A1_N(_05573_),
    .A2_N(_05589_),
    .B1(_05573_),
    .B2(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__nand2_2 _19897_ (.A(_05495_),
    .B(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__o21ai_2 _19898_ (.A1(_05495_),
    .A2(_05590_),
    .B1(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__or2_2 _19899_ (.A(_05564_),
    .B(_05592_),
    .X(_05593_));
 sky130_vsdinv _19900_ (.A(_05593_),
    .Y(_05594_));
 sky130_fd_sc_hd__a21o_2 _19901_ (.A1(_05564_),
    .A2(_05592_),
    .B1(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__o22a_2 _19902_ (.A1(_05539_),
    .A2(_05540_),
    .B1(_05525_),
    .B2(_05541_),
    .X(_05596_));
 sky130_fd_sc_hd__a21oi_2 _19903_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_05504_),
    .Y(_05597_));
 sky130_fd_sc_hd__buf_1 _19904_ (.A(_05508_),
    .X(_05598_));
 sky130_fd_sc_hd__buf_1 _19905_ (.A(_05598_),
    .X(_05599_));
 sky130_fd_sc_hd__o22a_2 _19906_ (.A1(_05153_),
    .A2(_05502_),
    .B1(_04694_),
    .B2(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__and4_2 _19907_ (.A(_11636_),
    .B(_11915_),
    .C(_11642_),
    .D(_11913_),
    .X(_05601_));
 sky130_fd_sc_hd__nor2_2 _19908_ (.A(_05600_),
    .B(_05601_),
    .Y(_05602_));
 sky130_fd_sc_hd__nor2_2 _19909_ (.A(_05251_),
    .B(_05421_),
    .Y(_05603_));
 sky130_fd_sc_hd__a2bb2o_2 _19910_ (.A1_N(_05602_),
    .A2_N(_05603_),
    .B1(_05602_),
    .B2(_05603_),
    .X(_05604_));
 sky130_vsdinv _19911_ (.A(\pcpi_mul.rs1[18] ),
    .Y(_05605_));
 sky130_fd_sc_hd__buf_1 _19912_ (.A(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__buf_1 _19913_ (.A(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__or2_2 _19914_ (.A(_04537_),
    .B(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__buf_1 _19915_ (.A(_05167_),
    .X(_05609_));
 sky130_fd_sc_hd__buf_1 _19916_ (.A(_05254_),
    .X(_05610_));
 sky130_fd_sc_hd__o22a_2 _19917_ (.A1(_05171_),
    .A2(_05609_),
    .B1(_05173_),
    .B2(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__buf_1 _19918_ (.A(\pcpi_mul.rs1[14] ),
    .X(_05612_));
 sky130_fd_sc_hd__and4_2 _19919_ (.A(_05513_),
    .B(_05516_),
    .C(_05515_),
    .D(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__or2_2 _19920_ (.A(_05611_),
    .B(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__a2bb2o_2 _19921_ (.A1_N(_05608_),
    .A2_N(_05614_),
    .B1(_05608_),
    .B2(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__o21ba_2 _19922_ (.A1(_05511_),
    .A2(_05518_),
    .B1_N(_05517_),
    .X(_05616_));
 sky130_fd_sc_hd__a2bb2o_2 _19923_ (.A1_N(_05615_),
    .A2_N(_05616_),
    .B1(_05615_),
    .B2(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__a2bb2o_2 _19924_ (.A1_N(_05604_),
    .A2_N(_05617_),
    .B1(_05604_),
    .B2(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__o22a_2 _19925_ (.A1(_05519_),
    .A2(_05520_),
    .B1(_05507_),
    .B2(_05521_),
    .X(_05619_));
 sky130_fd_sc_hd__a2bb2o_2 _19926_ (.A1_N(_05618_),
    .A2_N(_05619_),
    .B1(_05618_),
    .B2(_05619_),
    .X(_05620_));
 sky130_fd_sc_hd__a2bb2o_2 _19927_ (.A1_N(_05597_),
    .A2_N(_05620_),
    .B1(_05597_),
    .B2(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__o22a_2 _19928_ (.A1(_05529_),
    .A2(_05535_),
    .B1(_05528_),
    .B2(_05536_),
    .X(_05622_));
 sky130_fd_sc_hd__o22a_2 _19929_ (.A1(_05491_),
    .A2(_05492_),
    .B1(_05486_),
    .B2(_05493_),
    .X(_05623_));
 sky130_fd_sc_hd__o21ba_2 _19930_ (.A1(_05531_),
    .A2(_05534_),
    .B1_N(_05533_),
    .X(_05624_));
 sky130_fd_sc_hd__o21ba_2 _19931_ (.A1(_05482_),
    .A2(_05485_),
    .B1_N(_05484_),
    .X(_05625_));
 sky130_fd_sc_hd__or2_2 _19932_ (.A(_04829_),
    .B(_05157_),
    .X(_05626_));
 sky130_fd_sc_hd__o22a_2 _19933_ (.A1(_05275_),
    .A2(_05014_),
    .B1(_05276_),
    .B2(_05071_),
    .X(_05627_));
 sky130_fd_sc_hd__and4_2 _19934_ (.A(_05278_),
    .B(_11928_),
    .C(_05279_),
    .D(_11926_),
    .X(_05628_));
 sky130_fd_sc_hd__or2_2 _19935_ (.A(_05627_),
    .B(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__a2bb2o_2 _19936_ (.A1_N(_05626_),
    .A2_N(_05629_),
    .B1(_05626_),
    .B2(_05629_),
    .X(_05630_));
 sky130_fd_sc_hd__a2bb2o_2 _19937_ (.A1_N(_05625_),
    .A2_N(_05630_),
    .B1(_05625_),
    .B2(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__a2bb2o_2 _19938_ (.A1_N(_05624_),
    .A2_N(_05631_),
    .B1(_05624_),
    .B2(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__a2bb2o_2 _19939_ (.A1_N(_05623_),
    .A2_N(_05632_),
    .B1(_05623_),
    .B2(_05632_),
    .X(_05633_));
 sky130_fd_sc_hd__a2bb2o_2 _19940_ (.A1_N(_05622_),
    .A2_N(_05633_),
    .B1(_05622_),
    .B2(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__o22a_2 _19941_ (.A1(_05527_),
    .A2(_05537_),
    .B1(_05526_),
    .B2(_05538_),
    .X(_05635_));
 sky130_fd_sc_hd__a2bb2o_2 _19942_ (.A1_N(_05634_),
    .A2_N(_05635_),
    .B1(_05634_),
    .B2(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__a2bb2o_2 _19943_ (.A1_N(_05621_),
    .A2_N(_05636_),
    .B1(_05621_),
    .B2(_05636_),
    .X(_05637_));
 sky130_fd_sc_hd__a2bb2o_2 _19944_ (.A1_N(_05497_),
    .A2_N(_05637_),
    .B1(_05497_),
    .B2(_05637_),
    .X(_05638_));
 sky130_fd_sc_hd__a2bb2o_2 _19945_ (.A1_N(_05596_),
    .A2_N(_05638_),
    .B1(_05596_),
    .B2(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__or2_2 _19946_ (.A(_05595_),
    .B(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__a21bo_2 _19947_ (.A1(_05595_),
    .A2(_05639_),
    .B1_N(_05640_),
    .X(_05641_));
 sky130_fd_sc_hd__a2bb2o_2 _19948_ (.A1_N(_05545_),
    .A2_N(_05641_),
    .B1(_05545_),
    .B2(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__a2bb2o_2 _19949_ (.A1_N(_05559_),
    .A2_N(_05642_),
    .B1(_05559_),
    .B2(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__o22a_2 _19950_ (.A1(_05461_),
    .A2(_05546_),
    .B1(_05473_),
    .B2(_05547_),
    .X(_05644_));
 sky130_fd_sc_hd__a2bb2o_2 _19951_ (.A1_N(_05643_),
    .A2_N(_05644_),
    .B1(_05643_),
    .B2(_05644_),
    .X(_05645_));
 sky130_fd_sc_hd__a2bb2o_2 _19952_ (.A1_N(_05472_),
    .A2_N(_05645_),
    .B1(_05472_),
    .B2(_05645_),
    .X(_05646_));
 sky130_fd_sc_hd__o22a_2 _19953_ (.A1(_05548_),
    .A2(_05549_),
    .B1(_05385_),
    .B2(_05550_),
    .X(_05647_));
 sky130_fd_sc_hd__or2_2 _19954_ (.A(_05646_),
    .B(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__a21bo_2 _19955_ (.A1(_05646_),
    .A2(_05647_),
    .B1_N(_05648_),
    .X(_05649_));
 sky130_fd_sc_hd__a22o_2 _19956_ (.A1(_05551_),
    .A2(_05552_),
    .B1(_05469_),
    .B2(_05553_),
    .X(_05650_));
 sky130_fd_sc_hd__o31a_2 _19957_ (.A1(_05470_),
    .A2(_05554_),
    .A3(_05383_),
    .B1(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__a2bb2oi_2 _19958_ (.A1_N(_05649_),
    .A2_N(_05651_),
    .B1(_05649_),
    .B2(_05651_),
    .Y(_02637_));
 sky130_fd_sc_hd__o22a_2 _19959_ (.A1(_05643_),
    .A2(_05644_),
    .B1(_05472_),
    .B2(_05645_),
    .X(_05652_));
 sky130_fd_sc_hd__o22a_2 _19960_ (.A1(_05497_),
    .A2(_05637_),
    .B1(_05596_),
    .B2(_05638_),
    .X(_05653_));
 sky130_fd_sc_hd__o22a_2 _19961_ (.A1(_05618_),
    .A2(_05619_),
    .B1(_05597_),
    .B2(_05620_),
    .X(_05654_));
 sky130_fd_sc_hd__or2_2 _19962_ (.A(_05653_),
    .B(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__a21bo_2 _19963_ (.A1(_05653_),
    .A2(_05654_),
    .B1_N(_05655_),
    .X(_05656_));
 sky130_vsdinv _19964_ (.A(\pcpi_mul.rs2[19] ),
    .Y(_05657_));
 sky130_fd_sc_hd__buf_1 _19965_ (.A(_05657_),
    .X(_05658_));
 sky130_fd_sc_hd__buf_1 _19966_ (.A(_05658_),
    .X(_05659_));
 sky130_fd_sc_hd__buf_1 _19967_ (.A(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__o22a_2 _19968_ (.A1(_05660_),
    .A2(_04546_),
    .B1(_05563_),
    .B2(_04690_),
    .X(_05661_));
 sky130_fd_sc_hd__buf_1 _19969_ (.A(_05658_),
    .X(_05662_));
 sky130_fd_sc_hd__or4_2 _19970_ (.A(_05662_),
    .B(_04707_),
    .C(_05561_),
    .D(_04688_),
    .X(_05663_));
 sky130_fd_sc_hd__or2b_2 _19971_ (.A(_05661_),
    .B_N(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__buf_1 _19972_ (.A(_04953_),
    .X(_05665_));
 sky130_fd_sc_hd__or2_2 _19973_ (.A(_05665_),
    .B(_05070_),
    .X(_05666_));
 sky130_fd_sc_hd__buf_1 _19974_ (.A(_05140_),
    .X(_05667_));
 sky130_fd_sc_hd__o22a_2 _19975_ (.A1(_05060_),
    .A2(_05172_),
    .B1(_05667_),
    .B2(_05174_),
    .X(_05668_));
 sky130_fd_sc_hd__buf_1 _19976_ (.A(_05143_),
    .X(_05669_));
 sky130_fd_sc_hd__buf_1 _19977_ (.A(_11615_),
    .X(_05670_));
 sky130_fd_sc_hd__and4_2 _19978_ (.A(_05669_),
    .B(_05176_),
    .C(_05670_),
    .D(_05177_),
    .X(_05671_));
 sky130_fd_sc_hd__or2_2 _19979_ (.A(_05668_),
    .B(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__a2bb2o_2 _19980_ (.A1_N(_05666_),
    .A2_N(_05672_),
    .B1(_05666_),
    .B2(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__or2_2 _19981_ (.A(_05232_),
    .B(_05575_),
    .X(_05674_));
 sky130_fd_sc_hd__o22a_2 _19982_ (.A1(_05235_),
    .A2(_04876_),
    .B1(_05321_),
    .B2(_05100_),
    .X(_05675_));
 sky130_fd_sc_hd__and4_2 _19983_ (.A(_05323_),
    .B(_11942_),
    .C(_05237_),
    .D(_11938_),
    .X(_05676_));
 sky130_fd_sc_hd__or2_2 _19984_ (.A(_05675_),
    .B(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__a2bb2o_2 _19985_ (.A1_N(_05674_),
    .A2_N(_05677_),
    .B1(_05674_),
    .B2(_05677_),
    .X(_05678_));
 sky130_fd_sc_hd__o21ba_2 _19986_ (.A1(_05582_),
    .A2(_05585_),
    .B1_N(_05584_),
    .X(_05679_));
 sky130_fd_sc_hd__a2bb2o_2 _19987_ (.A1_N(_05678_),
    .A2_N(_05679_),
    .B1(_05678_),
    .B2(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__a2bb2o_2 _19988_ (.A1_N(_05673_),
    .A2_N(_05680_),
    .B1(_05673_),
    .B2(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__or2_2 _19989_ (.A(_05307_),
    .B(_04742_),
    .X(_05682_));
 sky130_fd_sc_hd__o22a_2 _19990_ (.A1(_05475_),
    .A2(_04699_),
    .B1(_05387_),
    .B2(_04721_),
    .X(_05683_));
 sky130_fd_sc_hd__and4_2 _19991_ (.A(_11601_),
    .B(_11950_),
    .C(\pcpi_mul.rs2[16] ),
    .D(_11947_),
    .X(_05684_));
 sky130_fd_sc_hd__or2_2 _19992_ (.A(_05683_),
    .B(_05684_),
    .X(_05685_));
 sky130_fd_sc_hd__a2bb2o_2 _19993_ (.A1_N(_05682_),
    .A2_N(_05685_),
    .B1(_05682_),
    .B2(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__o21ba_2 _19994_ (.A1(_05565_),
    .A2(_05568_),
    .B1_N(_05567_),
    .X(_05687_));
 sky130_fd_sc_hd__or2_2 _19995_ (.A(_05686_),
    .B(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__a21bo_2 _19996_ (.A1(_05686_),
    .A2(_05687_),
    .B1_N(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__a2bb2o_2 _19997_ (.A1_N(_05571_),
    .A2_N(_05689_),
    .B1(_05571_),
    .B2(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__a2bb2o_2 _19998_ (.A1_N(_05681_),
    .A2_N(_05690_),
    .B1(_05681_),
    .B2(_05690_),
    .X(_05691_));
 sky130_fd_sc_hd__o22a_2 _19999_ (.A1(_05480_),
    .A2(_05572_),
    .B1(_05573_),
    .B2(_05589_),
    .X(_05692_));
 sky130_fd_sc_hd__or2_2 _20000_ (.A(_05691_),
    .B(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__a21bo_2 _20001_ (.A1(_05691_),
    .A2(_05692_),
    .B1_N(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__or2_2 _20002_ (.A(_05664_),
    .B(_05694_),
    .X(_05695_));
 sky130_vsdinv _20003_ (.A(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__a21oi_2 _20004_ (.A1(_05664_),
    .A2(_05694_),
    .B1(_05696_),
    .Y(_05697_));
 sky130_vsdinv _20005_ (.A(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__a22o_2 _20006_ (.A1(_05593_),
    .A2(_05698_),
    .B1(_05594_),
    .B2(_05697_),
    .X(_05699_));
 sky130_fd_sc_hd__o22a_2 _20007_ (.A1(_05634_),
    .A2(_05635_),
    .B1(_05621_),
    .B2(_05636_),
    .X(_05700_));
 sky130_fd_sc_hd__a21oi_2 _20008_ (.A1(_05602_),
    .A2(_05603_),
    .B1(_05601_),
    .Y(_05701_));
 sky130_fd_sc_hd__buf_1 _20009_ (.A(_05153_),
    .X(_05702_));
 sky130_fd_sc_hd__buf_1 _20010_ (.A(_04694_),
    .X(_05703_));
 sky130_fd_sc_hd__buf_1 _20011_ (.A(_05607_),
    .X(_05704_));
 sky130_fd_sc_hd__o22a_2 _20012_ (.A1(_05702_),
    .A2(_05599_),
    .B1(_05703_),
    .B2(_05704_),
    .X(_05705_));
 sky130_fd_sc_hd__buf_1 _20013_ (.A(_11636_),
    .X(_05706_));
 sky130_fd_sc_hd__buf_1 _20014_ (.A(_11642_),
    .X(_05707_));
 sky130_fd_sc_hd__and4_2 _20015_ (.A(_05706_),
    .B(_11913_),
    .C(_05707_),
    .D(_11911_),
    .X(_05708_));
 sky130_fd_sc_hd__nor2_2 _20016_ (.A(_05705_),
    .B(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__buf_1 _20017_ (.A(_05251_),
    .X(_05710_));
 sky130_fd_sc_hd__nor2_2 _20018_ (.A(_05710_),
    .B(_05502_),
    .Y(_05711_));
 sky130_fd_sc_hd__a2bb2o_2 _20019_ (.A1_N(_05709_),
    .A2_N(_05711_),
    .B1(_05709_),
    .B2(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__buf_1 _20020_ (.A(_04719_),
    .X(_05713_));
 sky130_vsdinv _20021_ (.A(\pcpi_mul.rs1[19] ),
    .Y(_05714_));
 sky130_fd_sc_hd__buf_1 _20022_ (.A(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__buf_1 _20023_ (.A(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__or2_2 _20024_ (.A(_05713_),
    .B(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__buf_1 _20025_ (.A(_05171_),
    .X(_05718_));
 sky130_fd_sc_hd__buf_1 _20026_ (.A(_05173_),
    .X(_05719_));
 sky130_fd_sc_hd__buf_1 _20027_ (.A(_05342_),
    .X(_05720_));
 sky130_fd_sc_hd__o22a_2 _20028_ (.A1(_05718_),
    .A2(_05256_),
    .B1(_05719_),
    .B2(_05720_),
    .X(_05721_));
 sky130_fd_sc_hd__and4_2 _20029_ (.A(_11628_),
    .B(_11920_),
    .C(_11632_),
    .D(_11917_),
    .X(_05722_));
 sky130_fd_sc_hd__or2_2 _20030_ (.A(_05721_),
    .B(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__a2bb2o_2 _20031_ (.A1_N(_05717_),
    .A2_N(_05723_),
    .B1(_05717_),
    .B2(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__o21ba_2 _20032_ (.A1(_05608_),
    .A2(_05614_),
    .B1_N(_05613_),
    .X(_05725_));
 sky130_fd_sc_hd__a2bb2o_2 _20033_ (.A1_N(_05724_),
    .A2_N(_05725_),
    .B1(_05724_),
    .B2(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__a2bb2o_2 _20034_ (.A1_N(_05712_),
    .A2_N(_05726_),
    .B1(_05712_),
    .B2(_05726_),
    .X(_05727_));
 sky130_fd_sc_hd__o22a_2 _20035_ (.A1(_05615_),
    .A2(_05616_),
    .B1(_05604_),
    .B2(_05617_),
    .X(_05728_));
 sky130_fd_sc_hd__a2bb2o_2 _20036_ (.A1_N(_05727_),
    .A2_N(_05728_),
    .B1(_05727_),
    .B2(_05728_),
    .X(_05729_));
 sky130_fd_sc_hd__a2bb2o_2 _20037_ (.A1_N(_05701_),
    .A2_N(_05729_),
    .B1(_05701_),
    .B2(_05729_),
    .X(_05730_));
 sky130_fd_sc_hd__o22a_2 _20038_ (.A1(_05625_),
    .A2(_05630_),
    .B1(_05624_),
    .B2(_05631_),
    .X(_05731_));
 sky130_fd_sc_hd__o22a_2 _20039_ (.A1(_05586_),
    .A2(_05587_),
    .B1(_05581_),
    .B2(_05588_),
    .X(_05732_));
 sky130_fd_sc_hd__o21ba_2 _20040_ (.A1(_05626_),
    .A2(_05629_),
    .B1_N(_05628_),
    .X(_05733_));
 sky130_fd_sc_hd__o21ba_2 _20041_ (.A1(_05574_),
    .A2(_05580_),
    .B1_N(_05579_),
    .X(_05734_));
 sky130_fd_sc_hd__buf_1 _20042_ (.A(_04829_),
    .X(_05735_));
 sky130_fd_sc_hd__buf_1 _20043_ (.A(_05168_),
    .X(_05736_));
 sky130_fd_sc_hd__or2_2 _20044_ (.A(_05735_),
    .B(_05736_),
    .X(_05737_));
 sky130_fd_sc_hd__buf_1 _20045_ (.A(_05275_),
    .X(_05738_));
 sky130_fd_sc_hd__buf_1 _20046_ (.A(_05276_),
    .X(_05739_));
 sky130_fd_sc_hd__buf_1 _20047_ (.A(_05081_),
    .X(_05740_));
 sky130_fd_sc_hd__o22a_2 _20048_ (.A1(_05738_),
    .A2(_05154_),
    .B1(_05739_),
    .B2(_05740_),
    .X(_05741_));
 sky130_fd_sc_hd__buf_1 _20049_ (.A(_05278_),
    .X(_05742_));
 sky130_fd_sc_hd__buf_1 _20050_ (.A(\pcpi_mul.rs1[11] ),
    .X(_05743_));
 sky130_fd_sc_hd__buf_1 _20051_ (.A(_05279_),
    .X(_05744_));
 sky130_fd_sc_hd__buf_1 _20052_ (.A(\pcpi_mul.rs1[12] ),
    .X(_05745_));
 sky130_fd_sc_hd__and4_2 _20053_ (.A(_05742_),
    .B(_05743_),
    .C(_05744_),
    .D(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__or2_2 _20054_ (.A(_05741_),
    .B(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__a2bb2o_2 _20055_ (.A1_N(_05737_),
    .A2_N(_05747_),
    .B1(_05737_),
    .B2(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__a2bb2o_2 _20056_ (.A1_N(_05734_),
    .A2_N(_05748_),
    .B1(_05734_),
    .B2(_05748_),
    .X(_05749_));
 sky130_fd_sc_hd__a2bb2o_2 _20057_ (.A1_N(_05733_),
    .A2_N(_05749_),
    .B1(_05733_),
    .B2(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__a2bb2o_2 _20058_ (.A1_N(_05732_),
    .A2_N(_05750_),
    .B1(_05732_),
    .B2(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__a2bb2o_2 _20059_ (.A1_N(_05731_),
    .A2_N(_05751_),
    .B1(_05731_),
    .B2(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__o22a_2 _20060_ (.A1(_05623_),
    .A2(_05632_),
    .B1(_05622_),
    .B2(_05633_),
    .X(_05753_));
 sky130_fd_sc_hd__a2bb2o_2 _20061_ (.A1_N(_05752_),
    .A2_N(_05753_),
    .B1(_05752_),
    .B2(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__a2bb2o_2 _20062_ (.A1_N(_05730_),
    .A2_N(_05754_),
    .B1(_05730_),
    .B2(_05754_),
    .X(_05755_));
 sky130_fd_sc_hd__a2bb2o_2 _20063_ (.A1_N(_05591_),
    .A2_N(_05755_),
    .B1(_05591_),
    .B2(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__a2bb2o_2 _20064_ (.A1_N(_05700_),
    .A2_N(_05756_),
    .B1(_05700_),
    .B2(_05756_),
    .X(_05757_));
 sky130_fd_sc_hd__a2bb2o_2 _20065_ (.A1_N(_05699_),
    .A2_N(_05757_),
    .B1(_05699_),
    .B2(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__a2bb2o_2 _20066_ (.A1_N(_05640_),
    .A2_N(_05758_),
    .B1(_05640_),
    .B2(_05758_),
    .X(_05759_));
 sky130_fd_sc_hd__a2bb2o_2 _20067_ (.A1_N(_05656_),
    .A2_N(_05759_),
    .B1(_05656_),
    .B2(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__o22a_2 _20068_ (.A1(_05545_),
    .A2(_05641_),
    .B1(_05559_),
    .B2(_05642_),
    .X(_05761_));
 sky130_fd_sc_hd__a2bb2o_2 _20069_ (.A1_N(_05760_),
    .A2_N(_05761_),
    .B1(_05760_),
    .B2(_05761_),
    .X(_05762_));
 sky130_fd_sc_hd__a2bb2o_2 _20070_ (.A1_N(_05558_),
    .A2_N(_05762_),
    .B1(_05558_),
    .B2(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__and2_2 _20071_ (.A(_05652_),
    .B(_05763_),
    .X(_05764_));
 sky130_fd_sc_hd__or2_2 _20072_ (.A(_05652_),
    .B(_05763_),
    .X(_05765_));
 sky130_fd_sc_hd__or2b_2 _20073_ (.A(_05764_),
    .B_N(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__o21ai_2 _20074_ (.A1(_05649_),
    .A2(_05651_),
    .B1(_05648_),
    .Y(_05767_));
 sky130_fd_sc_hd__a2bb2o_2 _20075_ (.A1_N(_05766_),
    .A2_N(_05767_),
    .B1(_05766_),
    .B2(_05767_),
    .X(_02638_));
 sky130_fd_sc_hd__o22a_2 _20076_ (.A1(_05591_),
    .A2(_05755_),
    .B1(_05700_),
    .B2(_05756_),
    .X(_05768_));
 sky130_fd_sc_hd__o22a_2 _20077_ (.A1(_05727_),
    .A2(_05728_),
    .B1(_05701_),
    .B2(_05729_),
    .X(_05769_));
 sky130_fd_sc_hd__or2_2 _20078_ (.A(_05768_),
    .B(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__a21bo_2 _20079_ (.A1(_05768_),
    .A2(_05769_),
    .B1_N(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__or2_2 _20080_ (.A(_05560_),
    .B(_05061_),
    .X(_05772_));
 sky130_vsdinv _20081_ (.A(\pcpi_mul.rs2[20] ),
    .Y(_05773_));
 sky130_fd_sc_hd__o22a_2 _20082_ (.A1(_05657_),
    .A2(_04687_),
    .B1(_05773_),
    .B2(_04710_),
    .X(_05774_));
 sky130_fd_sc_hd__and4_2 _20083_ (.A(_11597_),
    .B(_11954_),
    .C(\pcpi_mul.rs2[20] ),
    .D(_11956_),
    .X(_05775_));
 sky130_fd_sc_hd__or2_2 _20084_ (.A(_05774_),
    .B(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__a2bb2o_2 _20085_ (.A1_N(_05772_),
    .A2_N(_05776_),
    .B1(_05772_),
    .B2(_05776_),
    .X(_05777_));
 sky130_fd_sc_hd__or2_2 _20086_ (.A(_05665_),
    .B(_05072_),
    .X(_05778_));
 sky130_fd_sc_hd__buf_1 _20087_ (.A(_05139_),
    .X(_05779_));
 sky130_fd_sc_hd__o22a_2 _20088_ (.A1(_05779_),
    .A2(_05174_),
    .B1(_05667_),
    .B2(_05258_),
    .X(_05780_));
 sky130_fd_sc_hd__buf_1 _20089_ (.A(_11930_),
    .X(_05781_));
 sky130_fd_sc_hd__and4_2 _20090_ (.A(_05669_),
    .B(_05781_),
    .C(_05670_),
    .D(_05260_),
    .X(_05782_));
 sky130_fd_sc_hd__or2_2 _20091_ (.A(_05780_),
    .B(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__a2bb2o_2 _20092_ (.A1_N(_05778_),
    .A2_N(_05783_),
    .B1(_05778_),
    .B2(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__or2_2 _20093_ (.A(_05056_),
    .B(_05017_),
    .X(_05785_));
 sky130_fd_sc_hd__o22a_2 _20094_ (.A1(_05405_),
    .A2(_05398_),
    .B1(_05131_),
    .B2(_05190_),
    .X(_05786_));
 sky130_fd_sc_hd__and4_2 _20095_ (.A(_11607_),
    .B(_11939_),
    .C(_11610_),
    .D(_05280_),
    .X(_05787_));
 sky130_fd_sc_hd__or2_2 _20096_ (.A(_05786_),
    .B(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__a2bb2o_2 _20097_ (.A1_N(_05785_),
    .A2_N(_05788_),
    .B1(_05785_),
    .B2(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__o21ba_2 _20098_ (.A1(_05674_),
    .A2(_05677_),
    .B1_N(_05676_),
    .X(_05790_));
 sky130_fd_sc_hd__a2bb2o_2 _20099_ (.A1_N(_05789_),
    .A2_N(_05790_),
    .B1(_05789_),
    .B2(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__a2bb2o_2 _20100_ (.A1_N(_05784_),
    .A2_N(_05791_),
    .B1(_05784_),
    .B2(_05791_),
    .X(_05792_));
 sky130_fd_sc_hd__o21ba_2 _20101_ (.A1(_05682_),
    .A2(_05685_),
    .B1_N(_05684_),
    .X(_05793_));
 sky130_fd_sc_hd__or2_2 _20102_ (.A(_05307_),
    .B(_05194_),
    .X(_05794_));
 sky130_fd_sc_hd__buf_1 _20103_ (.A(_05475_),
    .X(_05795_));
 sky130_fd_sc_hd__o22a_2 _20104_ (.A1(_05795_),
    .A2(_04782_),
    .B1(_05387_),
    .B2(_04742_),
    .X(_05796_));
 sky130_fd_sc_hd__and4_2 _20105_ (.A(_11601_),
    .B(_11948_),
    .C(_11604_),
    .D(_11945_),
    .X(_05797_));
 sky130_fd_sc_hd__or2_2 _20106_ (.A(_05796_),
    .B(_05797_),
    .X(_05798_));
 sky130_fd_sc_hd__a2bb2o_2 _20107_ (.A1_N(_05794_),
    .A2_N(_05798_),
    .B1(_05794_),
    .B2(_05798_),
    .X(_05799_));
 sky130_fd_sc_hd__a2bb2o_2 _20108_ (.A1_N(_05663_),
    .A2_N(_05799_),
    .B1(_05663_),
    .B2(_05799_),
    .X(_05800_));
 sky130_fd_sc_hd__a2bb2o_2 _20109_ (.A1_N(_05793_),
    .A2_N(_05800_),
    .B1(_05793_),
    .B2(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__a2bb2o_2 _20110_ (.A1_N(_05688_),
    .A2_N(_05801_),
    .B1(_05688_),
    .B2(_05801_),
    .X(_05802_));
 sky130_fd_sc_hd__a2bb2o_2 _20111_ (.A1_N(_05792_),
    .A2_N(_05802_),
    .B1(_05792_),
    .B2(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__o22a_2 _20112_ (.A1(_05571_),
    .A2(_05689_),
    .B1(_05681_),
    .B2(_05690_),
    .X(_05804_));
 sky130_fd_sc_hd__or2_2 _20113_ (.A(_05803_),
    .B(_05804_),
    .X(_05805_));
 sky130_fd_sc_hd__a21bo_2 _20114_ (.A1(_05803_),
    .A2(_05804_),
    .B1_N(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__or2_2 _20115_ (.A(_05777_),
    .B(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__a21bo_2 _20116_ (.A1(_05777_),
    .A2(_05806_),
    .B1_N(_05807_),
    .X(_05808_));
 sky130_vsdinv _20117_ (.A(_05808_),
    .Y(_05809_));
 sky130_fd_sc_hd__a22o_2 _20118_ (.A1(_05695_),
    .A2(_05808_),
    .B1(_05696_),
    .B2(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__o22a_2 _20119_ (.A1(_05752_),
    .A2(_05753_),
    .B1(_05730_),
    .B2(_05754_),
    .X(_05811_));
 sky130_fd_sc_hd__a21oi_2 _20120_ (.A1(_05709_),
    .A2(_05711_),
    .B1(_05708_),
    .Y(_05812_));
 sky130_fd_sc_hd__buf_1 _20121_ (.A(_05069_),
    .X(_05813_));
 sky130_fd_sc_hd__buf_1 _20122_ (.A(_05714_),
    .X(_05814_));
 sky130_fd_sc_hd__buf_1 _20123_ (.A(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__buf_1 _20124_ (.A(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__o22a_2 _20125_ (.A1(_05813_),
    .A2(_05704_),
    .B1(_05703_),
    .B2(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__and4_2 _20126_ (.A(_05706_),
    .B(_11911_),
    .C(_05707_),
    .D(_11909_),
    .X(_05818_));
 sky130_fd_sc_hd__nor2_2 _20127_ (.A(_05817_),
    .B(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__nor2_2 _20128_ (.A(_05710_),
    .B(_05599_),
    .Y(_05820_));
 sky130_fd_sc_hd__a2bb2o_2 _20129_ (.A1_N(_05819_),
    .A2_N(_05820_),
    .B1(_05819_),
    .B2(_05820_),
    .X(_05821_));
 sky130_vsdinv _20130_ (.A(\pcpi_mul.rs1[20] ),
    .Y(_05822_));
 sky130_fd_sc_hd__buf_1 _20131_ (.A(_05822_),
    .X(_05823_));
 sky130_fd_sc_hd__buf_1 _20132_ (.A(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__or2_2 _20133_ (.A(_04537_),
    .B(_05824_),
    .X(_05825_));
 sky130_fd_sc_hd__buf_1 _20134_ (.A(_05083_),
    .X(_05826_));
 sky130_fd_sc_hd__buf_1 _20135_ (.A(_05085_),
    .X(_05827_));
 sky130_fd_sc_hd__buf_1 _20136_ (.A(_05428_),
    .X(_05828_));
 sky130_fd_sc_hd__o22a_2 _20137_ (.A1(_05826_),
    .A2(_05343_),
    .B1(_05827_),
    .B2(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__buf_1 _20138_ (.A(\pcpi_mul.rs1[15] ),
    .X(_05830_));
 sky130_fd_sc_hd__buf_1 _20139_ (.A(_11914_),
    .X(_05831_));
 sky130_fd_sc_hd__and4_2 _20140_ (.A(_11628_),
    .B(_05830_),
    .C(_11632_),
    .D(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__or2_2 _20141_ (.A(_05829_),
    .B(_05832_),
    .X(_05833_));
 sky130_fd_sc_hd__a2bb2o_2 _20142_ (.A1_N(_05825_),
    .A2_N(_05833_),
    .B1(_05825_),
    .B2(_05833_),
    .X(_05834_));
 sky130_fd_sc_hd__o21ba_2 _20143_ (.A1(_05717_),
    .A2(_05723_),
    .B1_N(_05722_),
    .X(_05835_));
 sky130_fd_sc_hd__a2bb2o_2 _20144_ (.A1_N(_05834_),
    .A2_N(_05835_),
    .B1(_05834_),
    .B2(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__a2bb2o_2 _20145_ (.A1_N(_05821_),
    .A2_N(_05836_),
    .B1(_05821_),
    .B2(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__o22a_2 _20146_ (.A1(_05724_),
    .A2(_05725_),
    .B1(_05712_),
    .B2(_05726_),
    .X(_05838_));
 sky130_fd_sc_hd__a2bb2o_2 _20147_ (.A1_N(_05837_),
    .A2_N(_05838_),
    .B1(_05837_),
    .B2(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__a2bb2o_2 _20148_ (.A1_N(_05812_),
    .A2_N(_05839_),
    .B1(_05812_),
    .B2(_05839_),
    .X(_05840_));
 sky130_fd_sc_hd__o22a_2 _20149_ (.A1(_05734_),
    .A2(_05748_),
    .B1(_05733_),
    .B2(_05749_),
    .X(_05841_));
 sky130_fd_sc_hd__o22a_2 _20150_ (.A1(_05678_),
    .A2(_05679_),
    .B1(_05673_),
    .B2(_05680_),
    .X(_05842_));
 sky130_fd_sc_hd__o21ba_2 _20151_ (.A1(_05737_),
    .A2(_05747_),
    .B1_N(_05746_),
    .X(_05843_));
 sky130_fd_sc_hd__o21ba_2 _20152_ (.A1(_05666_),
    .A2(_05672_),
    .B1_N(_05671_),
    .X(_05844_));
 sky130_fd_sc_hd__buf_1 _20153_ (.A(_05610_),
    .X(_05845_));
 sky130_fd_sc_hd__or2_2 _20154_ (.A(_04794_),
    .B(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__o22a_2 _20155_ (.A1(_05193_),
    .A2(_05157_),
    .B1(_05739_),
    .B2(_05246_),
    .X(_05847_));
 sky130_fd_sc_hd__buf_1 _20156_ (.A(\pcpi_mul.rs1[13] ),
    .X(_05848_));
 sky130_fd_sc_hd__and4_2 _20157_ (.A(_05742_),
    .B(_05745_),
    .C(_05744_),
    .D(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__or2_2 _20158_ (.A(_05847_),
    .B(_05849_),
    .X(_05850_));
 sky130_fd_sc_hd__a2bb2o_2 _20159_ (.A1_N(_05846_),
    .A2_N(_05850_),
    .B1(_05846_),
    .B2(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__a2bb2o_2 _20160_ (.A1_N(_05844_),
    .A2_N(_05851_),
    .B1(_05844_),
    .B2(_05851_),
    .X(_05852_));
 sky130_fd_sc_hd__a2bb2o_2 _20161_ (.A1_N(_05843_),
    .A2_N(_05852_),
    .B1(_05843_),
    .B2(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__a2bb2o_2 _20162_ (.A1_N(_05842_),
    .A2_N(_05853_),
    .B1(_05842_),
    .B2(_05853_),
    .X(_05854_));
 sky130_fd_sc_hd__a2bb2o_2 _20163_ (.A1_N(_05841_),
    .A2_N(_05854_),
    .B1(_05841_),
    .B2(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__o22a_2 _20164_ (.A1(_05732_),
    .A2(_05750_),
    .B1(_05731_),
    .B2(_05751_),
    .X(_05856_));
 sky130_fd_sc_hd__a2bb2o_2 _20165_ (.A1_N(_05855_),
    .A2_N(_05856_),
    .B1(_05855_),
    .B2(_05856_),
    .X(_05857_));
 sky130_fd_sc_hd__a2bb2o_2 _20166_ (.A1_N(_05840_),
    .A2_N(_05857_),
    .B1(_05840_),
    .B2(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__a2bb2o_2 _20167_ (.A1_N(_05693_),
    .A2_N(_05858_),
    .B1(_05693_),
    .B2(_05858_),
    .X(_05859_));
 sky130_fd_sc_hd__a2bb2o_2 _20168_ (.A1_N(_05811_),
    .A2_N(_05859_),
    .B1(_05811_),
    .B2(_05859_),
    .X(_05860_));
 sky130_fd_sc_hd__a2bb2o_2 _20169_ (.A1_N(_05810_),
    .A2_N(_05860_),
    .B1(_05810_),
    .B2(_05860_),
    .X(_05861_));
 sky130_fd_sc_hd__o22a_2 _20170_ (.A1(_05593_),
    .A2(_05698_),
    .B1(_05699_),
    .B2(_05757_),
    .X(_05862_));
 sky130_fd_sc_hd__a2bb2o_2 _20171_ (.A1_N(_05861_),
    .A2_N(_05862_),
    .B1(_05861_),
    .B2(_05862_),
    .X(_05863_));
 sky130_fd_sc_hd__a2bb2o_2 _20172_ (.A1_N(_05771_),
    .A2_N(_05863_),
    .B1(_05771_),
    .B2(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__o22a_2 _20173_ (.A1(_05640_),
    .A2(_05758_),
    .B1(_05656_),
    .B2(_05759_),
    .X(_05865_));
 sky130_fd_sc_hd__a2bb2o_2 _20174_ (.A1_N(_05864_),
    .A2_N(_05865_),
    .B1(_05864_),
    .B2(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__a2bb2o_2 _20175_ (.A1_N(_05655_),
    .A2_N(_05866_),
    .B1(_05655_),
    .B2(_05866_),
    .X(_05867_));
 sky130_fd_sc_hd__o22a_2 _20176_ (.A1(_05760_),
    .A2(_05761_),
    .B1(_05558_),
    .B2(_05762_),
    .X(_05868_));
 sky130_fd_sc_hd__or2_2 _20177_ (.A(_05867_),
    .B(_05868_),
    .X(_05869_));
 sky130_fd_sc_hd__a21bo_2 _20178_ (.A1(_05867_),
    .A2(_05868_),
    .B1_N(_05869_),
    .X(_05870_));
 sky130_fd_sc_hd__or2_2 _20179_ (.A(_05649_),
    .B(_05766_),
    .X(_05871_));
 sky130_fd_sc_hd__or3_2 _20180_ (.A(_05470_),
    .B(_05554_),
    .C(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__o221a_2 _20181_ (.A1(_05648_),
    .A2(_05764_),
    .B1(_05650_),
    .B2(_05871_),
    .C1(_05765_),
    .X(_05873_));
 sky130_fd_sc_hd__o21ai_2 _20182_ (.A1(_05383_),
    .A2(_05872_),
    .B1(_05873_),
    .Y(_05874_));
 sky130_vsdinv _20183_ (.A(_05874_),
    .Y(_05875_));
 sky130_vsdinv _20184_ (.A(_05870_),
    .Y(_05876_));
 sky130_fd_sc_hd__o22a_2 _20185_ (.A1(_05870_),
    .A2(_05875_),
    .B1(_05876_),
    .B2(_05874_),
    .X(_02639_));
 sky130_fd_sc_hd__o22a_2 _20186_ (.A1(_05864_),
    .A2(_05865_),
    .B1(_05655_),
    .B2(_05866_),
    .X(_05877_));
 sky130_fd_sc_hd__o22a_2 _20187_ (.A1(_05693_),
    .A2(_05858_),
    .B1(_05811_),
    .B2(_05859_),
    .X(_05878_));
 sky130_fd_sc_hd__o22a_2 _20188_ (.A1(_05837_),
    .A2(_05838_),
    .B1(_05812_),
    .B2(_05839_),
    .X(_05879_));
 sky130_fd_sc_hd__or2_2 _20189_ (.A(_05878_),
    .B(_05879_),
    .X(_05880_));
 sky130_fd_sc_hd__a21bo_2 _20190_ (.A1(_05878_),
    .A2(_05879_),
    .B1_N(_05880_),
    .X(_05881_));
 sky130_fd_sc_hd__o22a_2 _20191_ (.A1(_05855_),
    .A2(_05856_),
    .B1(_05840_),
    .B2(_05857_),
    .X(_05882_));
 sky130_fd_sc_hd__a21oi_2 _20192_ (.A1(_05819_),
    .A2(_05820_),
    .B1(_05818_),
    .Y(_05883_));
 sky130_fd_sc_hd__buf_1 _20193_ (.A(_05822_),
    .X(_05884_));
 sky130_fd_sc_hd__buf_1 _20194_ (.A(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__o22a_2 _20195_ (.A1(_05813_),
    .A2(_05816_),
    .B1(_05703_),
    .B2(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__and4_2 _20196_ (.A(_05706_),
    .B(_11909_),
    .C(_05707_),
    .D(_11906_),
    .X(_05887_));
 sky130_fd_sc_hd__nor2_2 _20197_ (.A(_05886_),
    .B(_05887_),
    .Y(_05888_));
 sky130_fd_sc_hd__nor2_2 _20198_ (.A(_05710_),
    .B(_05704_),
    .Y(_05889_));
 sky130_fd_sc_hd__a2bb2o_2 _20199_ (.A1_N(_05888_),
    .A2_N(_05889_),
    .B1(_05888_),
    .B2(_05889_),
    .X(_05890_));
 sky130_vsdinv _20200_ (.A(\pcpi_mul.rs1[21] ),
    .Y(_05891_));
 sky130_fd_sc_hd__buf_1 _20201_ (.A(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__buf_1 _20202_ (.A(_05892_),
    .X(_05893_));
 sky130_fd_sc_hd__or2_2 _20203_ (.A(_04537_),
    .B(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__buf_1 _20204_ (.A(_05509_),
    .X(_05895_));
 sky130_fd_sc_hd__o22a_2 _20205_ (.A1(_05826_),
    .A2(_05429_),
    .B1(_05827_),
    .B2(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__buf_1 _20206_ (.A(\pcpi_mul.rs1[17] ),
    .X(_05897_));
 sky130_fd_sc_hd__and4_2 _20207_ (.A(_11628_),
    .B(_05831_),
    .C(_11632_),
    .D(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__or2_2 _20208_ (.A(_05896_),
    .B(_05898_),
    .X(_05899_));
 sky130_fd_sc_hd__a2bb2o_2 _20209_ (.A1_N(_05894_),
    .A2_N(_05899_),
    .B1(_05894_),
    .B2(_05899_),
    .X(_05900_));
 sky130_fd_sc_hd__o21ba_2 _20210_ (.A1(_05825_),
    .A2(_05833_),
    .B1_N(_05832_),
    .X(_05901_));
 sky130_fd_sc_hd__a2bb2o_2 _20211_ (.A1_N(_05900_),
    .A2_N(_05901_),
    .B1(_05900_),
    .B2(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__a2bb2o_2 _20212_ (.A1_N(_05890_),
    .A2_N(_05902_),
    .B1(_05890_),
    .B2(_05902_),
    .X(_05903_));
 sky130_fd_sc_hd__o22a_2 _20213_ (.A1(_05834_),
    .A2(_05835_),
    .B1(_05821_),
    .B2(_05836_),
    .X(_05904_));
 sky130_fd_sc_hd__a2bb2o_2 _20214_ (.A1_N(_05903_),
    .A2_N(_05904_),
    .B1(_05903_),
    .B2(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__a2bb2o_2 _20215_ (.A1_N(_05883_),
    .A2_N(_05905_),
    .B1(_05883_),
    .B2(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__o22a_2 _20216_ (.A1(_05844_),
    .A2(_05851_),
    .B1(_05843_),
    .B2(_05852_),
    .X(_05907_));
 sky130_fd_sc_hd__o22a_2 _20217_ (.A1(_05789_),
    .A2(_05790_),
    .B1(_05784_),
    .B2(_05791_),
    .X(_05908_));
 sky130_fd_sc_hd__o21ba_2 _20218_ (.A1(_05846_),
    .A2(_05850_),
    .B1_N(_05849_),
    .X(_05909_));
 sky130_fd_sc_hd__o21ba_2 _20219_ (.A1(_05778_),
    .A2(_05783_),
    .B1_N(_05782_),
    .X(_05910_));
 sky130_fd_sc_hd__or2_2 _20220_ (.A(_04794_),
    .B(_05720_),
    .X(_05911_));
 sky130_fd_sc_hd__o22a_2 _20221_ (.A1(_05193_),
    .A2(_05609_),
    .B1(_04827_),
    .B2(_05334_),
    .X(_05912_));
 sky130_fd_sc_hd__and4_2 _20222_ (.A(_11619_),
    .B(_05516_),
    .C(_11623_),
    .D(_05612_),
    .X(_05913_));
 sky130_fd_sc_hd__or2_2 _20223_ (.A(_05912_),
    .B(_05913_),
    .X(_05914_));
 sky130_fd_sc_hd__a2bb2o_2 _20224_ (.A1_N(_05911_),
    .A2_N(_05914_),
    .B1(_05911_),
    .B2(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__a2bb2o_2 _20225_ (.A1_N(_05910_),
    .A2_N(_05915_),
    .B1(_05910_),
    .B2(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__a2bb2o_2 _20226_ (.A1_N(_05909_),
    .A2_N(_05916_),
    .B1(_05909_),
    .B2(_05916_),
    .X(_05917_));
 sky130_fd_sc_hd__a2bb2o_2 _20227_ (.A1_N(_05908_),
    .A2_N(_05917_),
    .B1(_05908_),
    .B2(_05917_),
    .X(_05918_));
 sky130_fd_sc_hd__a2bb2o_2 _20228_ (.A1_N(_05907_),
    .A2_N(_05918_),
    .B1(_05907_),
    .B2(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__o22a_2 _20229_ (.A1(_05842_),
    .A2(_05853_),
    .B1(_05841_),
    .B2(_05854_),
    .X(_05920_));
 sky130_fd_sc_hd__a2bb2o_2 _20230_ (.A1_N(_05919_),
    .A2_N(_05920_),
    .B1(_05919_),
    .B2(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__a2bb2o_2 _20231_ (.A1_N(_05906_),
    .A2_N(_05921_),
    .B1(_05906_),
    .B2(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__a2bb2o_2 _20232_ (.A1_N(_05805_),
    .A2_N(_05922_),
    .B1(_05805_),
    .B2(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__a2bb2o_2 _20233_ (.A1_N(_05882_),
    .A2_N(_05923_),
    .B1(_05882_),
    .B2(_05923_),
    .X(_05924_));
 sky130_vsdinv _20234_ (.A(\pcpi_mul.rs2[21] ),
    .Y(_05925_));
 sky130_fd_sc_hd__buf_1 _20235_ (.A(_05925_),
    .X(_05926_));
 sky130_fd_sc_hd__buf_1 _20236_ (.A(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__or2_2 _20237_ (.A(_05927_),
    .B(_04544_),
    .X(_05928_));
 sky130_fd_sc_hd__or2_2 _20238_ (.A(_05560_),
    .B(_05406_),
    .X(_05929_));
 sky130_fd_sc_hd__o22a_2 _20239_ (.A1(_05773_),
    .A2(_04751_),
    .B1(_05657_),
    .B2(_04700_),
    .X(_05930_));
 sky130_fd_sc_hd__and4_2 _20240_ (.A(\pcpi_mul.rs2[20] ),
    .B(_05238_),
    .C(\pcpi_mul.rs2[19] ),
    .D(_11951_),
    .X(_05931_));
 sky130_fd_sc_hd__or2_2 _20241_ (.A(_05930_),
    .B(_05931_),
    .X(_05932_));
 sky130_fd_sc_hd__a2bb2o_2 _20242_ (.A1_N(_05929_),
    .A2_N(_05932_),
    .B1(_05929_),
    .B2(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__nor2_2 _20243_ (.A(_05928_),
    .B(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__a21o_2 _20244_ (.A1(_05928_),
    .A2(_05933_),
    .B1(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__o22a_2 _20245_ (.A1(_05688_),
    .A2(_05801_),
    .B1(_05792_),
    .B2(_05802_),
    .X(_05936_));
 sky130_fd_sc_hd__buf_1 _20246_ (.A(_05081_),
    .X(_05937_));
 sky130_fd_sc_hd__or2_2 _20247_ (.A(_05665_),
    .B(_05937_),
    .X(_05938_));
 sky130_fd_sc_hd__o22a_2 _20248_ (.A1(_05779_),
    .A2(_05163_),
    .B1(_05667_),
    .B2(_05154_),
    .X(_05939_));
 sky130_fd_sc_hd__and4_2 _20249_ (.A(_05669_),
    .B(_05260_),
    .C(_05670_),
    .D(_05433_),
    .X(_05940_));
 sky130_fd_sc_hd__or2_2 _20250_ (.A(_05939_),
    .B(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__a2bb2o_2 _20251_ (.A1_N(_05938_),
    .A2_N(_05941_),
    .B1(_05938_),
    .B2(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__buf_1 _20252_ (.A(_05013_),
    .X(_05943_));
 sky130_fd_sc_hd__or2_2 _20253_ (.A(_05133_),
    .B(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__buf_1 _20254_ (.A(_05234_),
    .X(_05945_));
 sky130_fd_sc_hd__o22a_2 _20255_ (.A1(_05945_),
    .A2(_05190_),
    .B1(_05131_),
    .B2(_05172_),
    .X(_05946_));
 sky130_fd_sc_hd__and4_2 _20256_ (.A(_11607_),
    .B(_05577_),
    .C(_11610_),
    .D(_05578_),
    .X(_05947_));
 sky130_fd_sc_hd__or2_2 _20257_ (.A(_05946_),
    .B(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__a2bb2o_2 _20258_ (.A1_N(_05944_),
    .A2_N(_05948_),
    .B1(_05944_),
    .B2(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__o21ba_2 _20259_ (.A1(_05785_),
    .A2(_05788_),
    .B1_N(_05787_),
    .X(_05950_));
 sky130_fd_sc_hd__a2bb2o_2 _20260_ (.A1_N(_05949_),
    .A2_N(_05950_),
    .B1(_05949_),
    .B2(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__a2bb2o_2 _20261_ (.A1_N(_05942_),
    .A2_N(_05951_),
    .B1(_05942_),
    .B2(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__o21ba_2 _20262_ (.A1(_05794_),
    .A2(_05798_),
    .B1_N(_05797_),
    .X(_05953_));
 sky130_fd_sc_hd__o21ba_2 _20263_ (.A1(_05772_),
    .A2(_05776_),
    .B1_N(_05775_),
    .X(_05954_));
 sky130_fd_sc_hd__or2_2 _20264_ (.A(_05308_),
    .B(_05195_),
    .X(_05955_));
 sky130_fd_sc_hd__o22a_2 _20265_ (.A1(_05795_),
    .A2(_04975_),
    .B1(_05391_),
    .B2(_05314_),
    .X(_05956_));
 sky130_fd_sc_hd__and4_2 _20266_ (.A(_11601_),
    .B(_11945_),
    .C(_11604_),
    .D(_11941_),
    .X(_05957_));
 sky130_fd_sc_hd__or2_2 _20267_ (.A(_05956_),
    .B(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__a2bb2o_2 _20268_ (.A1_N(_05955_),
    .A2_N(_05958_),
    .B1(_05955_),
    .B2(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__a2bb2o_2 _20269_ (.A1_N(_05954_),
    .A2_N(_05959_),
    .B1(_05954_),
    .B2(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__a2bb2o_2 _20270_ (.A1_N(_05953_),
    .A2_N(_05960_),
    .B1(_05953_),
    .B2(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__o22a_2 _20271_ (.A1(_05663_),
    .A2(_05799_),
    .B1(_05793_),
    .B2(_05800_),
    .X(_05962_));
 sky130_fd_sc_hd__a2bb2o_2 _20272_ (.A1_N(_05961_),
    .A2_N(_05962_),
    .B1(_05961_),
    .B2(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__a2bb2o_2 _20273_ (.A1_N(_05952_),
    .A2_N(_05963_),
    .B1(_05952_),
    .B2(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__or2_2 _20274_ (.A(_05936_),
    .B(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__a21bo_2 _20275_ (.A1(_05936_),
    .A2(_05964_),
    .B1_N(_05965_),
    .X(_05966_));
 sky130_fd_sc_hd__or2_2 _20276_ (.A(_05935_),
    .B(_05966_),
    .X(_05967_));
 sky130_fd_sc_hd__a21bo_2 _20277_ (.A1(_05935_),
    .A2(_05966_),
    .B1_N(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__a2bb2o_2 _20278_ (.A1_N(_05807_),
    .A2_N(_05968_),
    .B1(_05807_),
    .B2(_05968_),
    .X(_05969_));
 sky130_fd_sc_hd__a2bb2o_2 _20279_ (.A1_N(_05924_),
    .A2_N(_05969_),
    .B1(_05924_),
    .B2(_05969_),
    .X(_05970_));
 sky130_fd_sc_hd__o22a_2 _20280_ (.A1(_05695_),
    .A2(_05808_),
    .B1(_05810_),
    .B2(_05860_),
    .X(_05971_));
 sky130_fd_sc_hd__a2bb2o_2 _20281_ (.A1_N(_05970_),
    .A2_N(_05971_),
    .B1(_05970_),
    .B2(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__a2bb2o_2 _20282_ (.A1_N(_05881_),
    .A2_N(_05972_),
    .B1(_05881_),
    .B2(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__o22a_2 _20283_ (.A1(_05861_),
    .A2(_05862_),
    .B1(_05771_),
    .B2(_05863_),
    .X(_05974_));
 sky130_fd_sc_hd__a2bb2o_2 _20284_ (.A1_N(_05973_),
    .A2_N(_05974_),
    .B1(_05973_),
    .B2(_05974_),
    .X(_05975_));
 sky130_fd_sc_hd__a2bb2o_2 _20285_ (.A1_N(_05770_),
    .A2_N(_05975_),
    .B1(_05770_),
    .B2(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__or2_2 _20286_ (.A(_05877_),
    .B(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__a21bo_2 _20287_ (.A1(_05877_),
    .A2(_05976_),
    .B1_N(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__o21ai_2 _20288_ (.A1(_05870_),
    .A2(_05875_),
    .B1(_05869_),
    .Y(_05979_));
 sky130_fd_sc_hd__a2bb2o_2 _20289_ (.A1_N(_05978_),
    .A2_N(_05979_),
    .B1(_05978_),
    .B2(_05979_),
    .X(_02640_));
 sky130_fd_sc_hd__o22a_2 _20290_ (.A1(_05805_),
    .A2(_05922_),
    .B1(_05882_),
    .B2(_05923_),
    .X(_05980_));
 sky130_fd_sc_hd__o22a_2 _20291_ (.A1(_05903_),
    .A2(_05904_),
    .B1(_05883_),
    .B2(_05905_),
    .X(_05981_));
 sky130_fd_sc_hd__or2_2 _20292_ (.A(_05980_),
    .B(_05981_),
    .X(_05982_));
 sky130_fd_sc_hd__a21bo_2 _20293_ (.A1(_05980_),
    .A2(_05981_),
    .B1_N(_05982_),
    .X(_05983_));
 sky130_fd_sc_hd__o22a_2 _20294_ (.A1(_05919_),
    .A2(_05920_),
    .B1(_05906_),
    .B2(_05921_),
    .X(_05984_));
 sky130_fd_sc_hd__a21oi_2 _20295_ (.A1(_05888_),
    .A2(_05889_),
    .B1(_05887_),
    .Y(_05985_));
 sky130_fd_sc_hd__buf_1 _20296_ (.A(_05891_),
    .X(_05986_));
 sky130_fd_sc_hd__buf_1 _20297_ (.A(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__buf_1 _20298_ (.A(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__o22a_2 _20299_ (.A1(_05813_),
    .A2(_05885_),
    .B1(_05156_),
    .B2(_05988_),
    .X(_05989_));
 sky130_fd_sc_hd__and4_2 _20300_ (.A(_05706_),
    .B(_11906_),
    .C(_05707_),
    .D(_11903_),
    .X(_05990_));
 sky130_fd_sc_hd__nor2_2 _20301_ (.A(_05989_),
    .B(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__nor2_2 _20302_ (.A(_05710_),
    .B(_05816_),
    .Y(_05992_));
 sky130_fd_sc_hd__a2bb2o_2 _20303_ (.A1_N(_05991_),
    .A2_N(_05992_),
    .B1(_05991_),
    .B2(_05992_),
    .X(_05993_));
 sky130_vsdinv _20304_ (.A(\pcpi_mul.rs1[22] ),
    .Y(_05994_));
 sky130_fd_sc_hd__buf_1 _20305_ (.A(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__buf_1 _20306_ (.A(_05995_),
    .X(_05996_));
 sky130_fd_sc_hd__or2_2 _20307_ (.A(_04537_),
    .B(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__o22a_2 _20308_ (.A1(_05826_),
    .A2(_05895_),
    .B1(_05827_),
    .B2(_05607_),
    .X(_05998_));
 sky130_fd_sc_hd__buf_1 _20309_ (.A(\pcpi_mul.rs1[18] ),
    .X(_05999_));
 sky130_fd_sc_hd__and4_2 _20310_ (.A(_11628_),
    .B(_05897_),
    .C(_11632_),
    .D(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__or2_2 _20311_ (.A(_05998_),
    .B(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__a2bb2o_2 _20312_ (.A1_N(_05997_),
    .A2_N(_06001_),
    .B1(_05997_),
    .B2(_06001_),
    .X(_06002_));
 sky130_fd_sc_hd__o21ba_2 _20313_ (.A1(_05894_),
    .A2(_05899_),
    .B1_N(_05898_),
    .X(_06003_));
 sky130_fd_sc_hd__a2bb2o_2 _20314_ (.A1_N(_06002_),
    .A2_N(_06003_),
    .B1(_06002_),
    .B2(_06003_),
    .X(_06004_));
 sky130_fd_sc_hd__a2bb2o_2 _20315_ (.A1_N(_05993_),
    .A2_N(_06004_),
    .B1(_05993_),
    .B2(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__o22a_2 _20316_ (.A1(_05900_),
    .A2(_05901_),
    .B1(_05890_),
    .B2(_05902_),
    .X(_06006_));
 sky130_fd_sc_hd__a2bb2o_2 _20317_ (.A1_N(_06005_),
    .A2_N(_06006_),
    .B1(_06005_),
    .B2(_06006_),
    .X(_06007_));
 sky130_fd_sc_hd__a2bb2o_2 _20318_ (.A1_N(_05985_),
    .A2_N(_06007_),
    .B1(_05985_),
    .B2(_06007_),
    .X(_06008_));
 sky130_fd_sc_hd__o22a_2 _20319_ (.A1(_05910_),
    .A2(_05915_),
    .B1(_05909_),
    .B2(_05916_),
    .X(_06009_));
 sky130_fd_sc_hd__o22a_2 _20320_ (.A1(_05949_),
    .A2(_05950_),
    .B1(_05942_),
    .B2(_05951_),
    .X(_06010_));
 sky130_fd_sc_hd__o21ba_2 _20321_ (.A1(_05911_),
    .A2(_05914_),
    .B1_N(_05913_),
    .X(_06011_));
 sky130_fd_sc_hd__o21ba_2 _20322_ (.A1(_05938_),
    .A2(_05941_),
    .B1_N(_05940_),
    .X(_06012_));
 sky130_fd_sc_hd__or2_2 _20323_ (.A(_04794_),
    .B(_05828_),
    .X(_06013_));
 sky130_fd_sc_hd__buf_1 _20324_ (.A(_05341_),
    .X(_06014_));
 sky130_fd_sc_hd__o22a_2 _20325_ (.A1(_05193_),
    .A2(_05610_),
    .B1(_04827_),
    .B2(_06014_),
    .X(_06015_));
 sky130_fd_sc_hd__buf_1 _20326_ (.A(\pcpi_mul.rs1[15] ),
    .X(_06016_));
 sky130_fd_sc_hd__and4_2 _20327_ (.A(_11619_),
    .B(_05612_),
    .C(_11623_),
    .D(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__or2_2 _20328_ (.A(_06015_),
    .B(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__a2bb2o_2 _20329_ (.A1_N(_06013_),
    .A2_N(_06018_),
    .B1(_06013_),
    .B2(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__a2bb2o_2 _20330_ (.A1_N(_06012_),
    .A2_N(_06019_),
    .B1(_06012_),
    .B2(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__a2bb2o_2 _20331_ (.A1_N(_06011_),
    .A2_N(_06020_),
    .B1(_06011_),
    .B2(_06020_),
    .X(_06021_));
 sky130_fd_sc_hd__a2bb2o_2 _20332_ (.A1_N(_06010_),
    .A2_N(_06021_),
    .B1(_06010_),
    .B2(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__a2bb2o_2 _20333_ (.A1_N(_06009_),
    .A2_N(_06022_),
    .B1(_06009_),
    .B2(_06022_),
    .X(_06023_));
 sky130_fd_sc_hd__o22a_2 _20334_ (.A1(_05908_),
    .A2(_05917_),
    .B1(_05907_),
    .B2(_05918_),
    .X(_06024_));
 sky130_fd_sc_hd__a2bb2o_2 _20335_ (.A1_N(_06023_),
    .A2_N(_06024_),
    .B1(_06023_),
    .B2(_06024_),
    .X(_06025_));
 sky130_fd_sc_hd__a2bb2o_2 _20336_ (.A1_N(_06008_),
    .A2_N(_06025_),
    .B1(_06008_),
    .B2(_06025_),
    .X(_06026_));
 sky130_fd_sc_hd__a2bb2o_2 _20337_ (.A1_N(_05965_),
    .A2_N(_06026_),
    .B1(_05965_),
    .B2(_06026_),
    .X(_06027_));
 sky130_fd_sc_hd__a2bb2o_2 _20338_ (.A1_N(_05984_),
    .A2_N(_06027_),
    .B1(_05984_),
    .B2(_06027_),
    .X(_06028_));
 sky130_vsdinv _20339_ (.A(\pcpi_mul.rs2[22] ),
    .Y(_06029_));
 sky130_fd_sc_hd__buf_1 _20340_ (.A(_06029_),
    .X(_06030_));
 sky130_fd_sc_hd__buf_1 _20341_ (.A(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__o22a_2 _20342_ (.A1(_06031_),
    .A2(_04543_),
    .B1(_05926_),
    .B2(_04689_),
    .X(_06032_));
 sky130_fd_sc_hd__buf_1 _20343_ (.A(_06029_),
    .X(_06033_));
 sky130_fd_sc_hd__buf_1 _20344_ (.A(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__buf_1 _20345_ (.A(_05925_),
    .X(_06035_));
 sky130_fd_sc_hd__or4_2 _20346_ (.A(_06034_),
    .B(_04707_),
    .C(_06035_),
    .D(_04703_),
    .X(_06036_));
 sky130_fd_sc_hd__or2b_2 _20347_ (.A(_06032_),
    .B_N(_06036_),
    .X(_06037_));
 sky130_fd_sc_hd__or2_2 _20348_ (.A(_05561_),
    .B(_05403_),
    .X(_06038_));
 sky130_fd_sc_hd__buf_1 _20349_ (.A(_05773_),
    .X(_06039_));
 sky130_fd_sc_hd__o22a_2 _20350_ (.A1(_06039_),
    .A2(_04779_),
    .B1(_05658_),
    .B2(_05141_),
    .X(_06040_));
 sky130_fd_sc_hd__and4_2 _20351_ (.A(_11592_),
    .B(_05144_),
    .C(_11597_),
    .D(_05145_),
    .X(_06041_));
 sky130_fd_sc_hd__or2_2 _20352_ (.A(_06040_),
    .B(_06041_),
    .X(_06042_));
 sky130_fd_sc_hd__a2bb2o_2 _20353_ (.A1_N(_06038_),
    .A2_N(_06042_),
    .B1(_06038_),
    .B2(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__or2_2 _20354_ (.A(_06037_),
    .B(_06043_),
    .X(_06044_));
 sky130_fd_sc_hd__a21boi_2 _20355_ (.A1(_06037_),
    .A2(_06043_),
    .B1_N(_06044_),
    .Y(_06045_));
 sky130_fd_sc_hd__nand2_2 _20356_ (.A(_05934_),
    .B(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__o21ai_2 _20357_ (.A1(_05934_),
    .A2(_06045_),
    .B1(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__o22a_2 _20358_ (.A1(_05961_),
    .A2(_05962_),
    .B1(_05952_),
    .B2(_05963_),
    .X(_06048_));
 sky130_fd_sc_hd__buf_1 _20359_ (.A(_04902_),
    .X(_06049_));
 sky130_fd_sc_hd__or2_2 _20360_ (.A(_06049_),
    .B(_05247_),
    .X(_06050_));
 sky130_fd_sc_hd__buf_1 _20361_ (.A(_05060_),
    .X(_06051_));
 sky130_fd_sc_hd__buf_1 _20362_ (.A(_04950_),
    .X(_06052_));
 sky130_fd_sc_hd__o22a_2 _20363_ (.A1(_06051_),
    .A2(_05154_),
    .B1(_06052_),
    .B2(_05740_),
    .X(_06053_));
 sky130_fd_sc_hd__buf_1 _20364_ (.A(_11613_),
    .X(_06054_));
 sky130_fd_sc_hd__buf_1 _20365_ (.A(_11616_),
    .X(_06055_));
 sky130_fd_sc_hd__and4_2 _20366_ (.A(_06054_),
    .B(_05743_),
    .C(_06055_),
    .D(_05745_),
    .X(_06056_));
 sky130_fd_sc_hd__or2_2 _20367_ (.A(_06053_),
    .B(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__a2bb2o_2 _20368_ (.A1_N(_06050_),
    .A2_N(_06057_),
    .B1(_06050_),
    .B2(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__or2_2 _20369_ (.A(_05133_),
    .B(_05070_),
    .X(_06059_));
 sky130_fd_sc_hd__o22a_2 _20370_ (.A1(_05945_),
    .A2(_05172_),
    .B1(_05131_),
    .B2(_05076_),
    .X(_06060_));
 sky130_fd_sc_hd__and4_2 _20371_ (.A(_11607_),
    .B(_05578_),
    .C(_11610_),
    .D(_05177_),
    .X(_06061_));
 sky130_fd_sc_hd__or2_2 _20372_ (.A(_06060_),
    .B(_06061_),
    .X(_06062_));
 sky130_fd_sc_hd__a2bb2o_2 _20373_ (.A1_N(_06059_),
    .A2_N(_06062_),
    .B1(_06059_),
    .B2(_06062_),
    .X(_06063_));
 sky130_fd_sc_hd__o21ba_2 _20374_ (.A1(_05944_),
    .A2(_05948_),
    .B1_N(_05947_),
    .X(_06064_));
 sky130_fd_sc_hd__a2bb2o_2 _20375_ (.A1_N(_06063_),
    .A2_N(_06064_),
    .B1(_06063_),
    .B2(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__a2bb2o_2 _20376_ (.A1_N(_06058_),
    .A2_N(_06065_),
    .B1(_06058_),
    .B2(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__o21ba_2 _20377_ (.A1(_05955_),
    .A2(_05958_),
    .B1_N(_05957_),
    .X(_06067_));
 sky130_fd_sc_hd__o21ba_2 _20378_ (.A1(_05929_),
    .A2(_05932_),
    .B1_N(_05931_),
    .X(_06068_));
 sky130_fd_sc_hd__or2_2 _20379_ (.A(_05308_),
    .B(_05575_),
    .X(_06069_));
 sky130_fd_sc_hd__o22a_2 _20380_ (.A1(_05795_),
    .A2(_04876_),
    .B1(_05391_),
    .B2(_05100_),
    .X(_06070_));
 sky130_fd_sc_hd__and4_2 _20381_ (.A(_11601_),
    .B(_11942_),
    .C(_11604_),
    .D(_11938_),
    .X(_06071_));
 sky130_fd_sc_hd__or2_2 _20382_ (.A(_06070_),
    .B(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__a2bb2o_2 _20383_ (.A1_N(_06069_),
    .A2_N(_06072_),
    .B1(_06069_),
    .B2(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__a2bb2o_2 _20384_ (.A1_N(_06068_),
    .A2_N(_06073_),
    .B1(_06068_),
    .B2(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__a2bb2o_2 _20385_ (.A1_N(_06067_),
    .A2_N(_06074_),
    .B1(_06067_),
    .B2(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__o22a_2 _20386_ (.A1(_05954_),
    .A2(_05959_),
    .B1(_05953_),
    .B2(_05960_),
    .X(_06076_));
 sky130_fd_sc_hd__a2bb2o_2 _20387_ (.A1_N(_06075_),
    .A2_N(_06076_),
    .B1(_06075_),
    .B2(_06076_),
    .X(_06077_));
 sky130_fd_sc_hd__a2bb2o_2 _20388_ (.A1_N(_06066_),
    .A2_N(_06077_),
    .B1(_06066_),
    .B2(_06077_),
    .X(_06078_));
 sky130_fd_sc_hd__or2_2 _20389_ (.A(_06048_),
    .B(_06078_),
    .X(_06079_));
 sky130_fd_sc_hd__a21bo_2 _20390_ (.A1(_06048_),
    .A2(_06078_),
    .B1_N(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__or2_2 _20391_ (.A(_06047_),
    .B(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__a21bo_2 _20392_ (.A1(_06047_),
    .A2(_06080_),
    .B1_N(_06081_),
    .X(_06082_));
 sky130_fd_sc_hd__a2bb2o_2 _20393_ (.A1_N(_05967_),
    .A2_N(_06082_),
    .B1(_05967_),
    .B2(_06082_),
    .X(_06083_));
 sky130_fd_sc_hd__a2bb2o_2 _20394_ (.A1_N(_06028_),
    .A2_N(_06083_),
    .B1(_06028_),
    .B2(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__o22a_2 _20395_ (.A1(_05807_),
    .A2(_05968_),
    .B1(_05924_),
    .B2(_05969_),
    .X(_06085_));
 sky130_fd_sc_hd__a2bb2o_2 _20396_ (.A1_N(_06084_),
    .A2_N(_06085_),
    .B1(_06084_),
    .B2(_06085_),
    .X(_06086_));
 sky130_fd_sc_hd__a2bb2o_2 _20397_ (.A1_N(_05983_),
    .A2_N(_06086_),
    .B1(_05983_),
    .B2(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__o22a_2 _20398_ (.A1(_05970_),
    .A2(_05971_),
    .B1(_05881_),
    .B2(_05972_),
    .X(_06088_));
 sky130_fd_sc_hd__a2bb2o_2 _20399_ (.A1_N(_06087_),
    .A2_N(_06088_),
    .B1(_06087_),
    .B2(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__a2bb2o_2 _20400_ (.A1_N(_05880_),
    .A2_N(_06089_),
    .B1(_05880_),
    .B2(_06089_),
    .X(_06090_));
 sky130_fd_sc_hd__o22a_2 _20401_ (.A1(_05973_),
    .A2(_05974_),
    .B1(_05770_),
    .B2(_05975_),
    .X(_06091_));
 sky130_fd_sc_hd__or2_2 _20402_ (.A(_06090_),
    .B(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__a21bo_2 _20403_ (.A1(_06090_),
    .A2(_06091_),
    .B1_N(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__a22o_2 _20404_ (.A1(_05877_),
    .A2(_05976_),
    .B1(_05869_),
    .B2(_05977_),
    .X(_06094_));
 sky130_fd_sc_hd__o31a_2 _20405_ (.A1(_05870_),
    .A2(_05978_),
    .A3(_05875_),
    .B1(_06094_),
    .X(_06095_));
 sky130_fd_sc_hd__a2bb2oi_2 _20406_ (.A1_N(_06093_),
    .A2_N(_06095_),
    .B1(_06093_),
    .B2(_06095_),
    .Y(_02641_));
 sky130_fd_sc_hd__o22a_2 _20407_ (.A1(_06087_),
    .A2(_06088_),
    .B1(_05880_),
    .B2(_06089_),
    .X(_06096_));
 sky130_fd_sc_hd__o22a_2 _20408_ (.A1(_05965_),
    .A2(_06026_),
    .B1(_05984_),
    .B2(_06027_),
    .X(_06097_));
 sky130_fd_sc_hd__o22a_2 _20409_ (.A1(_06005_),
    .A2(_06006_),
    .B1(_05985_),
    .B2(_06007_),
    .X(_06098_));
 sky130_fd_sc_hd__or2_2 _20410_ (.A(_06097_),
    .B(_06098_),
    .X(_06099_));
 sky130_fd_sc_hd__a21bo_2 _20411_ (.A1(_06097_),
    .A2(_06098_),
    .B1_N(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__o22a_2 _20412_ (.A1(_06023_),
    .A2(_06024_),
    .B1(_06008_),
    .B2(_06025_),
    .X(_06101_));
 sky130_fd_sc_hd__a21oi_2 _20413_ (.A1(_05991_),
    .A2(_05992_),
    .B1(_05990_),
    .Y(_06102_));
 sky130_fd_sc_hd__buf_1 _20414_ (.A(_05996_),
    .X(_06103_));
 sky130_fd_sc_hd__o22a_2 _20415_ (.A1(_05702_),
    .A2(_05988_),
    .B1(_04695_),
    .B2(_06103_),
    .X(_06104_));
 sky130_fd_sc_hd__and4_2 _20416_ (.A(_11638_),
    .B(_11903_),
    .C(_11644_),
    .D(_11901_),
    .X(_06105_));
 sky130_fd_sc_hd__nor2_2 _20417_ (.A(_06104_),
    .B(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__buf_1 _20418_ (.A(_05162_),
    .X(_06107_));
 sky130_fd_sc_hd__nor2_2 _20419_ (.A(_06107_),
    .B(_05885_),
    .Y(_06108_));
 sky130_fd_sc_hd__a2bb2o_2 _20420_ (.A1_N(_06106_),
    .A2_N(_06108_),
    .B1(_06106_),
    .B2(_06108_),
    .X(_06109_));
 sky130_vsdinv _20421_ (.A(\pcpi_mul.rs1[23] ),
    .Y(_06110_));
 sky130_fd_sc_hd__buf_1 _20422_ (.A(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__buf_1 _20423_ (.A(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__or2_2 _20424_ (.A(_04538_),
    .B(_06112_),
    .X(_06113_));
 sky130_fd_sc_hd__o22a_2 _20425_ (.A1(_05718_),
    .A2(_05607_),
    .B1(_05719_),
    .B2(_05815_),
    .X(_06114_));
 sky130_fd_sc_hd__buf_1 _20426_ (.A(_05513_),
    .X(_06115_));
 sky130_fd_sc_hd__buf_1 _20427_ (.A(_05515_),
    .X(_06116_));
 sky130_fd_sc_hd__buf_1 _20428_ (.A(\pcpi_mul.rs1[19] ),
    .X(_06117_));
 sky130_fd_sc_hd__and4_2 _20429_ (.A(_06115_),
    .B(_11911_),
    .C(_06116_),
    .D(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__or2_2 _20430_ (.A(_06114_),
    .B(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__a2bb2o_2 _20431_ (.A1_N(_06113_),
    .A2_N(_06119_),
    .B1(_06113_),
    .B2(_06119_),
    .X(_06120_));
 sky130_fd_sc_hd__o21ba_2 _20432_ (.A1(_05997_),
    .A2(_06001_),
    .B1_N(_06000_),
    .X(_06121_));
 sky130_fd_sc_hd__a2bb2o_2 _20433_ (.A1_N(_06120_),
    .A2_N(_06121_),
    .B1(_06120_),
    .B2(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__a2bb2o_2 _20434_ (.A1_N(_06109_),
    .A2_N(_06122_),
    .B1(_06109_),
    .B2(_06122_),
    .X(_06123_));
 sky130_fd_sc_hd__o22a_2 _20435_ (.A1(_06002_),
    .A2(_06003_),
    .B1(_05993_),
    .B2(_06004_),
    .X(_06124_));
 sky130_fd_sc_hd__a2bb2o_2 _20436_ (.A1_N(_06123_),
    .A2_N(_06124_),
    .B1(_06123_),
    .B2(_06124_),
    .X(_06125_));
 sky130_fd_sc_hd__a2bb2o_2 _20437_ (.A1_N(_06102_),
    .A2_N(_06125_),
    .B1(_06102_),
    .B2(_06125_),
    .X(_06126_));
 sky130_fd_sc_hd__o22a_2 _20438_ (.A1(_06012_),
    .A2(_06019_),
    .B1(_06011_),
    .B2(_06020_),
    .X(_06127_));
 sky130_fd_sc_hd__o22a_2 _20439_ (.A1(_06063_),
    .A2(_06064_),
    .B1(_06058_),
    .B2(_06065_),
    .X(_06128_));
 sky130_fd_sc_hd__o21ba_2 _20440_ (.A1(_06013_),
    .A2(_06018_),
    .B1_N(_06017_),
    .X(_06129_));
 sky130_fd_sc_hd__o21ba_2 _20441_ (.A1(_06050_),
    .A2(_06057_),
    .B1_N(_06056_),
    .X(_06130_));
 sky130_fd_sc_hd__or2_2 _20442_ (.A(_04830_),
    .B(_05510_),
    .X(_06131_));
 sky130_fd_sc_hd__buf_1 _20443_ (.A(_05275_),
    .X(_06132_));
 sky130_fd_sc_hd__buf_1 _20444_ (.A(_05276_),
    .X(_06133_));
 sky130_fd_sc_hd__buf_1 _20445_ (.A(_05428_),
    .X(_06134_));
 sky130_fd_sc_hd__o22a_2 _20446_ (.A1(_06132_),
    .A2(_06014_),
    .B1(_06133_),
    .B2(_06134_),
    .X(_06135_));
 sky130_fd_sc_hd__buf_1 _20447_ (.A(_11619_),
    .X(_06136_));
 sky130_fd_sc_hd__buf_1 _20448_ (.A(_11623_),
    .X(_06137_));
 sky130_fd_sc_hd__buf_1 _20449_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06138_));
 sky130_fd_sc_hd__and4_2 _20450_ (.A(_06136_),
    .B(_06016_),
    .C(_06137_),
    .D(_06138_),
    .X(_06139_));
 sky130_fd_sc_hd__or2_2 _20451_ (.A(_06135_),
    .B(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__a2bb2o_2 _20452_ (.A1_N(_06131_),
    .A2_N(_06140_),
    .B1(_06131_),
    .B2(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__a2bb2o_2 _20453_ (.A1_N(_06130_),
    .A2_N(_06141_),
    .B1(_06130_),
    .B2(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__a2bb2o_2 _20454_ (.A1_N(_06129_),
    .A2_N(_06142_),
    .B1(_06129_),
    .B2(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__a2bb2o_2 _20455_ (.A1_N(_06128_),
    .A2_N(_06143_),
    .B1(_06128_),
    .B2(_06143_),
    .X(_06144_));
 sky130_fd_sc_hd__a2bb2o_2 _20456_ (.A1_N(_06127_),
    .A2_N(_06144_),
    .B1(_06127_),
    .B2(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__o22a_2 _20457_ (.A1(_06010_),
    .A2(_06021_),
    .B1(_06009_),
    .B2(_06022_),
    .X(_06146_));
 sky130_fd_sc_hd__a2bb2o_2 _20458_ (.A1_N(_06145_),
    .A2_N(_06146_),
    .B1(_06145_),
    .B2(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__a2bb2o_2 _20459_ (.A1_N(_06126_),
    .A2_N(_06147_),
    .B1(_06126_),
    .B2(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__a2bb2o_2 _20460_ (.A1_N(_06079_),
    .A2_N(_06148_),
    .B1(_06079_),
    .B2(_06148_),
    .X(_06149_));
 sky130_fd_sc_hd__a2bb2o_2 _20461_ (.A1_N(_06101_),
    .A2_N(_06149_),
    .B1(_06101_),
    .B2(_06149_),
    .X(_06150_));
 sky130_fd_sc_hd__buf_1 _20462_ (.A(_05314_),
    .X(_06151_));
 sky130_fd_sc_hd__or2_2 _20463_ (.A(_05561_),
    .B(_06151_),
    .X(_06152_));
 sky130_fd_sc_hd__o22a_2 _20464_ (.A1(_06039_),
    .A2(_05141_),
    .B1(_05658_),
    .B2(_05227_),
    .X(_06153_));
 sky130_fd_sc_hd__and4_2 _20465_ (.A(_11592_),
    .B(_11949_),
    .C(_11597_),
    .D(_05316_),
    .X(_06154_));
 sky130_fd_sc_hd__or2_2 _20466_ (.A(_06153_),
    .B(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__a2bb2o_2 _20467_ (.A1_N(_06152_),
    .A2_N(_06155_),
    .B1(_06152_),
    .B2(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__or2_2 _20468_ (.A(_05925_),
    .B(_04702_),
    .X(_06157_));
 sky130_vsdinv _20469_ (.A(\pcpi_mul.rs2[23] ),
    .Y(_06158_));
 sky130_fd_sc_hd__o22a_2 _20470_ (.A1(_06029_),
    .A2(_04751_),
    .B1(_06158_),
    .B2(_04710_),
    .X(_06159_));
 sky130_fd_sc_hd__and4_2 _20471_ (.A(_11588_),
    .B(_05238_),
    .C(\pcpi_mul.rs2[23] ),
    .D(_11957_),
    .X(_06160_));
 sky130_fd_sc_hd__or2_2 _20472_ (.A(_06159_),
    .B(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__a2bb2o_2 _20473_ (.A1_N(_06157_),
    .A2_N(_06161_),
    .B1(_06157_),
    .B2(_06161_),
    .X(_06162_));
 sky130_fd_sc_hd__a2bb2o_2 _20474_ (.A1_N(_06036_),
    .A2_N(_06162_),
    .B1(_06036_),
    .B2(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__a2bb2o_2 _20475_ (.A1_N(_06156_),
    .A2_N(_06163_),
    .B1(_06156_),
    .B2(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__or2_2 _20476_ (.A(_06044_),
    .B(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__a21bo_2 _20477_ (.A1(_06044_),
    .A2(_06164_),
    .B1_N(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__o22a_2 _20478_ (.A1(_06075_),
    .A2(_06076_),
    .B1(_06066_),
    .B2(_06077_),
    .X(_06167_));
 sky130_fd_sc_hd__buf_1 _20479_ (.A(_04902_),
    .X(_06168_));
 sky130_fd_sc_hd__or2_2 _20480_ (.A(_06168_),
    .B(_05845_),
    .X(_06169_));
 sky130_fd_sc_hd__o22a_2 _20481_ (.A1(_06051_),
    .A2(_05431_),
    .B1(_06052_),
    .B2(_05246_),
    .X(_06170_));
 sky130_fd_sc_hd__buf_1 _20482_ (.A(_11613_),
    .X(_06171_));
 sky130_fd_sc_hd__buf_1 _20483_ (.A(_11616_),
    .X(_06172_));
 sky130_fd_sc_hd__and4_2 _20484_ (.A(_06171_),
    .B(_05514_),
    .C(_06172_),
    .D(_05516_),
    .X(_06173_));
 sky130_fd_sc_hd__or2_2 _20485_ (.A(_06170_),
    .B(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__a2bb2o_2 _20486_ (.A1_N(_06169_),
    .A2_N(_06174_),
    .B1(_06169_),
    .B2(_06174_),
    .X(_06175_));
 sky130_fd_sc_hd__buf_1 _20487_ (.A(_05232_),
    .X(_06176_));
 sky130_fd_sc_hd__or2_2 _20488_ (.A(_06176_),
    .B(_05072_),
    .X(_06177_));
 sky130_fd_sc_hd__buf_1 _20489_ (.A(_05405_),
    .X(_06178_));
 sky130_fd_sc_hd__buf_1 _20490_ (.A(_05321_),
    .X(_06179_));
 sky130_fd_sc_hd__buf_1 _20491_ (.A(_05014_),
    .X(_06180_));
 sky130_fd_sc_hd__o22a_2 _20492_ (.A1(_06178_),
    .A2(_05174_),
    .B1(_06179_),
    .B2(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__buf_1 _20493_ (.A(_05323_),
    .X(_06182_));
 sky130_fd_sc_hd__buf_1 _20494_ (.A(_05237_),
    .X(_06183_));
 sky130_fd_sc_hd__buf_1 _20495_ (.A(_11928_),
    .X(_06184_));
 sky130_fd_sc_hd__and4_2 _20496_ (.A(_06182_),
    .B(_05781_),
    .C(_06183_),
    .D(_06184_),
    .X(_06185_));
 sky130_fd_sc_hd__or2_2 _20497_ (.A(_06181_),
    .B(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__a2bb2o_2 _20498_ (.A1_N(_06177_),
    .A2_N(_06186_),
    .B1(_06177_),
    .B2(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__o21ba_2 _20499_ (.A1(_06059_),
    .A2(_06062_),
    .B1_N(_06061_),
    .X(_06188_));
 sky130_fd_sc_hd__a2bb2o_2 _20500_ (.A1_N(_06187_),
    .A2_N(_06188_),
    .B1(_06187_),
    .B2(_06188_),
    .X(_06189_));
 sky130_fd_sc_hd__a2bb2o_2 _20501_ (.A1_N(_06175_),
    .A2_N(_06189_),
    .B1(_06175_),
    .B2(_06189_),
    .X(_06190_));
 sky130_fd_sc_hd__o21ba_2 _20502_ (.A1(_06069_),
    .A2(_06072_),
    .B1_N(_06071_),
    .X(_06191_));
 sky130_fd_sc_hd__o21ba_2 _20503_ (.A1(_06038_),
    .A2(_06042_),
    .B1_N(_06041_),
    .X(_06192_));
 sky130_fd_sc_hd__or2_2 _20504_ (.A(_05308_),
    .B(_05017_),
    .X(_06193_));
 sky130_fd_sc_hd__o22a_2 _20505_ (.A1(_05795_),
    .A2(_05398_),
    .B1(_05391_),
    .B2(_05084_),
    .X(_06194_));
 sky130_fd_sc_hd__and4_2 _20506_ (.A(_11602_),
    .B(_11939_),
    .C(_11605_),
    .D(_05280_),
    .X(_06195_));
 sky130_fd_sc_hd__or2_2 _20507_ (.A(_06194_),
    .B(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__a2bb2o_2 _20508_ (.A1_N(_06193_),
    .A2_N(_06196_),
    .B1(_06193_),
    .B2(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__a2bb2o_2 _20509_ (.A1_N(_06192_),
    .A2_N(_06197_),
    .B1(_06192_),
    .B2(_06197_),
    .X(_06198_));
 sky130_fd_sc_hd__a2bb2o_2 _20510_ (.A1_N(_06191_),
    .A2_N(_06198_),
    .B1(_06191_),
    .B2(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__o22a_2 _20511_ (.A1(_06068_),
    .A2(_06073_),
    .B1(_06067_),
    .B2(_06074_),
    .X(_06200_));
 sky130_fd_sc_hd__a2bb2o_2 _20512_ (.A1_N(_06199_),
    .A2_N(_06200_),
    .B1(_06199_),
    .B2(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__a2bb2o_2 _20513_ (.A1_N(_06190_),
    .A2_N(_06201_),
    .B1(_06190_),
    .B2(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__a2bb2o_2 _20514_ (.A1_N(_06046_),
    .A2_N(_06202_),
    .B1(_06046_),
    .B2(_06202_),
    .X(_06203_));
 sky130_fd_sc_hd__a2bb2o_2 _20515_ (.A1_N(_06167_),
    .A2_N(_06203_),
    .B1(_06167_),
    .B2(_06203_),
    .X(_06204_));
 sky130_fd_sc_hd__or2_2 _20516_ (.A(_06166_),
    .B(_06204_),
    .X(_06205_));
 sky130_fd_sc_hd__a21bo_2 _20517_ (.A1(_06166_),
    .A2(_06204_),
    .B1_N(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__a2bb2o_2 _20518_ (.A1_N(_06081_),
    .A2_N(_06206_),
    .B1(_06081_),
    .B2(_06206_),
    .X(_06207_));
 sky130_fd_sc_hd__a2bb2o_2 _20519_ (.A1_N(_06150_),
    .A2_N(_06207_),
    .B1(_06150_),
    .B2(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__o22a_2 _20520_ (.A1(_05967_),
    .A2(_06082_),
    .B1(_06028_),
    .B2(_06083_),
    .X(_06209_));
 sky130_fd_sc_hd__a2bb2o_2 _20521_ (.A1_N(_06208_),
    .A2_N(_06209_),
    .B1(_06208_),
    .B2(_06209_),
    .X(_06210_));
 sky130_fd_sc_hd__a2bb2o_2 _20522_ (.A1_N(_06100_),
    .A2_N(_06210_),
    .B1(_06100_),
    .B2(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__o22a_2 _20523_ (.A1(_06084_),
    .A2(_06085_),
    .B1(_05983_),
    .B2(_06086_),
    .X(_06212_));
 sky130_fd_sc_hd__a2bb2o_2 _20524_ (.A1_N(_06211_),
    .A2_N(_06212_),
    .B1(_06211_),
    .B2(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__a2bb2o_2 _20525_ (.A1_N(_05982_),
    .A2_N(_06213_),
    .B1(_05982_),
    .B2(_06213_),
    .X(_06214_));
 sky130_fd_sc_hd__and2_2 _20526_ (.A(_06096_),
    .B(_06214_),
    .X(_06215_));
 sky130_fd_sc_hd__or2_2 _20527_ (.A(_06096_),
    .B(_06214_),
    .X(_06216_));
 sky130_fd_sc_hd__or2b_2 _20528_ (.A(_06215_),
    .B_N(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__o21ai_2 _20529_ (.A1(_06093_),
    .A2(_06095_),
    .B1(_06092_),
    .Y(_06218_));
 sky130_fd_sc_hd__a2bb2o_2 _20530_ (.A1_N(_06217_),
    .A2_N(_06218_),
    .B1(_06217_),
    .B2(_06218_),
    .X(_02642_));
 sky130_fd_sc_hd__o22a_2 _20531_ (.A1(_06079_),
    .A2(_06148_),
    .B1(_06101_),
    .B2(_06149_),
    .X(_06219_));
 sky130_fd_sc_hd__o22a_2 _20532_ (.A1(_06123_),
    .A2(_06124_),
    .B1(_06102_),
    .B2(_06125_),
    .X(_06220_));
 sky130_fd_sc_hd__or2_2 _20533_ (.A(_06219_),
    .B(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__a21bo_2 _20534_ (.A1(_06219_),
    .A2(_06220_),
    .B1_N(_06221_),
    .X(_06222_));
 sky130_fd_sc_hd__o22a_2 _20535_ (.A1(_06145_),
    .A2(_06146_),
    .B1(_06126_),
    .B2(_06147_),
    .X(_06223_));
 sky130_fd_sc_hd__o22a_2 _20536_ (.A1(_06046_),
    .A2(_06202_),
    .B1(_06167_),
    .B2(_06203_),
    .X(_06224_));
 sky130_fd_sc_hd__a21oi_2 _20537_ (.A1(_06106_),
    .A2(_06108_),
    .B1(_06105_),
    .Y(_06225_));
 sky130_fd_sc_hd__buf_1 _20538_ (.A(_06112_),
    .X(_06226_));
 sky130_fd_sc_hd__o22a_2 _20539_ (.A1(_05702_),
    .A2(_06103_),
    .B1(_04695_),
    .B2(_06226_),
    .X(_06227_));
 sky130_fd_sc_hd__and4_2 _20540_ (.A(_11638_),
    .B(_11901_),
    .C(_11644_),
    .D(_11898_),
    .X(_06228_));
 sky130_fd_sc_hd__nor2_2 _20541_ (.A(_06227_),
    .B(_06228_),
    .Y(_06229_));
 sky130_fd_sc_hd__nor2_2 _20542_ (.A(_06107_),
    .B(_05988_),
    .Y(_06230_));
 sky130_fd_sc_hd__a2bb2o_2 _20543_ (.A1_N(_06229_),
    .A2_N(_06230_),
    .B1(_06229_),
    .B2(_06230_),
    .X(_06231_));
 sky130_vsdinv _20544_ (.A(\pcpi_mul.rs1[24] ),
    .Y(_06232_));
 sky130_fd_sc_hd__buf_1 _20545_ (.A(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__buf_1 _20546_ (.A(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__or2_2 _20547_ (.A(_05713_),
    .B(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__buf_1 _20548_ (.A(_05822_),
    .X(_06236_));
 sky130_fd_sc_hd__buf_1 _20549_ (.A(_06236_),
    .X(_06237_));
 sky130_fd_sc_hd__o22a_2 _20550_ (.A1(_05718_),
    .A2(_05815_),
    .B1(_05719_),
    .B2(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__buf_1 _20551_ (.A(\pcpi_mul.rs1[20] ),
    .X(_06239_));
 sky130_fd_sc_hd__buf_1 _20552_ (.A(_06239_),
    .X(_06240_));
 sky130_fd_sc_hd__and4_2 _20553_ (.A(_06115_),
    .B(_06117_),
    .C(_06116_),
    .D(_06240_),
    .X(_06241_));
 sky130_fd_sc_hd__or2_2 _20554_ (.A(_06238_),
    .B(_06241_),
    .X(_06242_));
 sky130_fd_sc_hd__a2bb2o_2 _20555_ (.A1_N(_06235_),
    .A2_N(_06242_),
    .B1(_06235_),
    .B2(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__o21ba_2 _20556_ (.A1(_06113_),
    .A2(_06119_),
    .B1_N(_06118_),
    .X(_06244_));
 sky130_fd_sc_hd__a2bb2o_2 _20557_ (.A1_N(_06243_),
    .A2_N(_06244_),
    .B1(_06243_),
    .B2(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__a2bb2o_2 _20558_ (.A1_N(_06231_),
    .A2_N(_06245_),
    .B1(_06231_),
    .B2(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__o22a_2 _20559_ (.A1(_06120_),
    .A2(_06121_),
    .B1(_06109_),
    .B2(_06122_),
    .X(_06247_));
 sky130_fd_sc_hd__a2bb2o_2 _20560_ (.A1_N(_06246_),
    .A2_N(_06247_),
    .B1(_06246_),
    .B2(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__a2bb2o_2 _20561_ (.A1_N(_06225_),
    .A2_N(_06248_),
    .B1(_06225_),
    .B2(_06248_),
    .X(_06249_));
 sky130_fd_sc_hd__o22a_2 _20562_ (.A1(_06130_),
    .A2(_06141_),
    .B1(_06129_),
    .B2(_06142_),
    .X(_06250_));
 sky130_fd_sc_hd__o22a_2 _20563_ (.A1(_06187_),
    .A2(_06188_),
    .B1(_06175_),
    .B2(_06189_),
    .X(_06251_));
 sky130_fd_sc_hd__o21ba_2 _20564_ (.A1(_06131_),
    .A2(_06140_),
    .B1_N(_06139_),
    .X(_06252_));
 sky130_fd_sc_hd__o21ba_2 _20565_ (.A1(_06169_),
    .A2(_06174_),
    .B1_N(_06173_),
    .X(_06253_));
 sky130_fd_sc_hd__buf_1 _20566_ (.A(_05605_),
    .X(_06254_));
 sky130_fd_sc_hd__buf_1 _20567_ (.A(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__or2_2 _20568_ (.A(_05735_),
    .B(_06255_),
    .X(_06256_));
 sky130_fd_sc_hd__buf_1 _20569_ (.A(_05508_),
    .X(_06257_));
 sky130_fd_sc_hd__o22a_2 _20570_ (.A1(_05738_),
    .A2(_05501_),
    .B1(_06133_),
    .B2(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__and4_2 _20571_ (.A(_05742_),
    .B(_06138_),
    .C(_05744_),
    .D(_11912_),
    .X(_06259_));
 sky130_fd_sc_hd__or2_2 _20572_ (.A(_06258_),
    .B(_06259_),
    .X(_06260_));
 sky130_fd_sc_hd__a2bb2o_2 _20573_ (.A1_N(_06256_),
    .A2_N(_06260_),
    .B1(_06256_),
    .B2(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__a2bb2o_2 _20574_ (.A1_N(_06253_),
    .A2_N(_06261_),
    .B1(_06253_),
    .B2(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__a2bb2o_2 _20575_ (.A1_N(_06252_),
    .A2_N(_06262_),
    .B1(_06252_),
    .B2(_06262_),
    .X(_06263_));
 sky130_fd_sc_hd__a2bb2o_2 _20576_ (.A1_N(_06251_),
    .A2_N(_06263_),
    .B1(_06251_),
    .B2(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__a2bb2o_2 _20577_ (.A1_N(_06250_),
    .A2_N(_06264_),
    .B1(_06250_),
    .B2(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__o22a_2 _20578_ (.A1(_06128_),
    .A2(_06143_),
    .B1(_06127_),
    .B2(_06144_),
    .X(_06266_));
 sky130_fd_sc_hd__a2bb2o_2 _20579_ (.A1_N(_06265_),
    .A2_N(_06266_),
    .B1(_06265_),
    .B2(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__a2bb2o_2 _20580_ (.A1_N(_06249_),
    .A2_N(_06267_),
    .B1(_06249_),
    .B2(_06267_),
    .X(_06268_));
 sky130_fd_sc_hd__a2bb2o_2 _20581_ (.A1_N(_06224_),
    .A2_N(_06268_),
    .B1(_06224_),
    .B2(_06268_),
    .X(_06269_));
 sky130_fd_sc_hd__a2bb2o_2 _20582_ (.A1_N(_06223_),
    .A2_N(_06269_),
    .B1(_06223_),
    .B2(_06269_),
    .X(_06270_));
 sky130_vsdinv _20583_ (.A(\pcpi_mul.rs2[24] ),
    .Y(_06271_));
 sky130_fd_sc_hd__buf_1 _20584_ (.A(_06271_),
    .X(_06272_));
 sky130_fd_sc_hd__buf_1 _20585_ (.A(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__buf_1 _20586_ (.A(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__buf_1 _20587_ (.A(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__or2_2 _20588_ (.A(_06275_),
    .B(_04545_),
    .X(_06276_));
 sky130_fd_sc_hd__buf_1 _20589_ (.A(_05398_),
    .X(_06277_));
 sky130_fd_sc_hd__or2_2 _20590_ (.A(_05561_),
    .B(_06277_),
    .X(_06278_));
 sky130_fd_sc_hd__o22a_2 _20591_ (.A1(_06039_),
    .A2(_05137_),
    .B1(_05658_),
    .B2(_05225_),
    .X(_06279_));
 sky130_fd_sc_hd__buf_1 _20592_ (.A(_11597_),
    .X(_06280_));
 sky130_fd_sc_hd__and4_2 _20593_ (.A(_11592_),
    .B(_11946_),
    .C(_06280_),
    .D(_05197_),
    .X(_06281_));
 sky130_fd_sc_hd__or2_2 _20594_ (.A(_06279_),
    .B(_06281_),
    .X(_06282_));
 sky130_fd_sc_hd__a2bb2o_2 _20595_ (.A1_N(_06278_),
    .A2_N(_06282_),
    .B1(_06278_),
    .B2(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__or2_2 _20596_ (.A(_05925_),
    .B(_05406_),
    .X(_06284_));
 sky130_fd_sc_hd__o22a_2 _20597_ (.A1(_06158_),
    .A2(_04751_),
    .B1(_06029_),
    .B2(_04701_),
    .X(_06285_));
 sky130_fd_sc_hd__and4_2 _20598_ (.A(\pcpi_mul.rs2[23] ),
    .B(_05238_),
    .C(\pcpi_mul.rs2[22] ),
    .D(_11951_),
    .X(_06286_));
 sky130_fd_sc_hd__or2_2 _20599_ (.A(_06285_),
    .B(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__a2bb2o_2 _20600_ (.A1_N(_06284_),
    .A2_N(_06287_),
    .B1(_06284_),
    .B2(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__o21ba_2 _20601_ (.A1(_06157_),
    .A2(_06161_),
    .B1_N(_06160_),
    .X(_06289_));
 sky130_fd_sc_hd__a2bb2o_2 _20602_ (.A1_N(_06288_),
    .A2_N(_06289_),
    .B1(_06288_),
    .B2(_06289_),
    .X(_06290_));
 sky130_fd_sc_hd__a2bb2o_2 _20603_ (.A1_N(_06283_),
    .A2_N(_06290_),
    .B1(_06283_),
    .B2(_06290_),
    .X(_06291_));
 sky130_fd_sc_hd__o22a_2 _20604_ (.A1(_06036_),
    .A2(_06162_),
    .B1(_06156_),
    .B2(_06163_),
    .X(_06292_));
 sky130_fd_sc_hd__or2_2 _20605_ (.A(_06291_),
    .B(_06292_),
    .X(_06293_));
 sky130_fd_sc_hd__a21bo_2 _20606_ (.A1(_06291_),
    .A2(_06292_),
    .B1_N(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__or2_2 _20607_ (.A(_06276_),
    .B(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__a21bo_2 _20608_ (.A1(_06276_),
    .A2(_06294_),
    .B1_N(_06295_),
    .X(_06296_));
 sky130_fd_sc_hd__o22a_2 _20609_ (.A1(_06199_),
    .A2(_06200_),
    .B1(_06190_),
    .B2(_06201_),
    .X(_06297_));
 sky130_fd_sc_hd__or2_2 _20610_ (.A(_06168_),
    .B(_05720_),
    .X(_06298_));
 sky130_fd_sc_hd__buf_1 _20611_ (.A(_05139_),
    .X(_06299_));
 sky130_fd_sc_hd__buf_1 _20612_ (.A(_05140_),
    .X(_06300_));
 sky130_fd_sc_hd__o22a_2 _20613_ (.A1(_06299_),
    .A2(_05609_),
    .B1(_06300_),
    .B2(_05610_),
    .X(_06301_));
 sky130_fd_sc_hd__and4_2 _20614_ (.A(_06171_),
    .B(_05516_),
    .C(_06172_),
    .D(_05612_),
    .X(_06302_));
 sky130_fd_sc_hd__or2_2 _20615_ (.A(_06301_),
    .B(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__a2bb2o_2 _20616_ (.A1_N(_06298_),
    .A2_N(_06303_),
    .B1(_06298_),
    .B2(_06303_),
    .X(_06304_));
 sky130_fd_sc_hd__buf_1 _20617_ (.A(_05056_),
    .X(_06305_));
 sky130_fd_sc_hd__or2_2 _20618_ (.A(_06305_),
    .B(_05937_),
    .X(_06306_));
 sky130_fd_sc_hd__buf_1 _20619_ (.A(_05235_),
    .X(_06307_));
 sky130_fd_sc_hd__o22a_2 _20620_ (.A1(_06307_),
    .A2(_05258_),
    .B1(_06179_),
    .B2(_05154_),
    .X(_06308_));
 sky130_fd_sc_hd__and4_2 _20621_ (.A(_06182_),
    .B(_06184_),
    .C(_06183_),
    .D(_05433_),
    .X(_06309_));
 sky130_fd_sc_hd__or2_2 _20622_ (.A(_06308_),
    .B(_06309_),
    .X(_06310_));
 sky130_fd_sc_hd__a2bb2o_2 _20623_ (.A1_N(_06306_),
    .A2_N(_06310_),
    .B1(_06306_),
    .B2(_06310_),
    .X(_06311_));
 sky130_fd_sc_hd__o21ba_2 _20624_ (.A1(_06177_),
    .A2(_06186_),
    .B1_N(_06185_),
    .X(_06312_));
 sky130_fd_sc_hd__a2bb2o_2 _20625_ (.A1_N(_06311_),
    .A2_N(_06312_),
    .B1(_06311_),
    .B2(_06312_),
    .X(_06313_));
 sky130_fd_sc_hd__a2bb2o_2 _20626_ (.A1_N(_06304_),
    .A2_N(_06313_),
    .B1(_06304_),
    .B2(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__o21ba_2 _20627_ (.A1(_06193_),
    .A2(_06196_),
    .B1_N(_06195_),
    .X(_06315_));
 sky130_fd_sc_hd__o21ba_2 _20628_ (.A1(_06152_),
    .A2(_06155_),
    .B1_N(_06154_),
    .X(_06316_));
 sky130_fd_sc_hd__or2_2 _20629_ (.A(_05308_),
    .B(_05943_),
    .X(_06317_));
 sky130_fd_sc_hd__buf_1 _20630_ (.A(_05795_),
    .X(_06318_));
 sky130_fd_sc_hd__o22a_2 _20631_ (.A1(_06318_),
    .A2(_05190_),
    .B1(_05391_),
    .B2(_05086_),
    .X(_06319_));
 sky130_fd_sc_hd__and4_2 _20632_ (.A(_11602_),
    .B(_05280_),
    .C(_11605_),
    .D(_05578_),
    .X(_06320_));
 sky130_fd_sc_hd__or2_2 _20633_ (.A(_06319_),
    .B(_06320_),
    .X(_06321_));
 sky130_fd_sc_hd__a2bb2o_2 _20634_ (.A1_N(_06317_),
    .A2_N(_06321_),
    .B1(_06317_),
    .B2(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__a2bb2o_2 _20635_ (.A1_N(_06316_),
    .A2_N(_06322_),
    .B1(_06316_),
    .B2(_06322_),
    .X(_06323_));
 sky130_fd_sc_hd__a2bb2o_2 _20636_ (.A1_N(_06315_),
    .A2_N(_06323_),
    .B1(_06315_),
    .B2(_06323_),
    .X(_06324_));
 sky130_fd_sc_hd__o22a_2 _20637_ (.A1(_06192_),
    .A2(_06197_),
    .B1(_06191_),
    .B2(_06198_),
    .X(_06325_));
 sky130_fd_sc_hd__a2bb2o_2 _20638_ (.A1_N(_06324_),
    .A2_N(_06325_),
    .B1(_06324_),
    .B2(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__a2bb2o_2 _20639_ (.A1_N(_06314_),
    .A2_N(_06326_),
    .B1(_06314_),
    .B2(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__a2bb2o_2 _20640_ (.A1_N(_06165_),
    .A2_N(_06327_),
    .B1(_06165_),
    .B2(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__a2bb2o_2 _20641_ (.A1_N(_06297_),
    .A2_N(_06328_),
    .B1(_06297_),
    .B2(_06328_),
    .X(_06329_));
 sky130_fd_sc_hd__or2_2 _20642_ (.A(_06296_),
    .B(_06329_),
    .X(_06330_));
 sky130_fd_sc_hd__a21bo_2 _20643_ (.A1(_06296_),
    .A2(_06329_),
    .B1_N(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__a2bb2o_2 _20644_ (.A1_N(_06205_),
    .A2_N(_06331_),
    .B1(_06205_),
    .B2(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__a2bb2o_2 _20645_ (.A1_N(_06270_),
    .A2_N(_06332_),
    .B1(_06270_),
    .B2(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__o22a_2 _20646_ (.A1(_06081_),
    .A2(_06206_),
    .B1(_06150_),
    .B2(_06207_),
    .X(_06334_));
 sky130_fd_sc_hd__a2bb2o_2 _20647_ (.A1_N(_06333_),
    .A2_N(_06334_),
    .B1(_06333_),
    .B2(_06334_),
    .X(_06335_));
 sky130_fd_sc_hd__a2bb2o_2 _20648_ (.A1_N(_06222_),
    .A2_N(_06335_),
    .B1(_06222_),
    .B2(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__o22a_2 _20649_ (.A1(_06208_),
    .A2(_06209_),
    .B1(_06100_),
    .B2(_06210_),
    .X(_06337_));
 sky130_fd_sc_hd__a2bb2o_2 _20650_ (.A1_N(_06336_),
    .A2_N(_06337_),
    .B1(_06336_),
    .B2(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__a2bb2o_2 _20651_ (.A1_N(_06099_),
    .A2_N(_06338_),
    .B1(_06099_),
    .B2(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__o22a_2 _20652_ (.A1(_06211_),
    .A2(_06212_),
    .B1(_05982_),
    .B2(_06213_),
    .X(_06340_));
 sky130_fd_sc_hd__or2_2 _20653_ (.A(_06339_),
    .B(_06340_),
    .X(_06341_));
 sky130_fd_sc_hd__a21bo_2 _20654_ (.A1(_06339_),
    .A2(_06340_),
    .B1_N(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__or2_2 _20655_ (.A(_06093_),
    .B(_06217_),
    .X(_06343_));
 sky130_fd_sc_hd__or3_2 _20656_ (.A(_05870_),
    .B(_05978_),
    .C(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__or3_2 _20657_ (.A(_05872_),
    .B(_06344_),
    .C(_05383_),
    .X(_06345_));
 sky130_fd_sc_hd__o21a_2 _20658_ (.A1(_06092_),
    .A2(_06215_),
    .B1(_06216_),
    .X(_06346_));
 sky130_fd_sc_hd__o221a_2 _20659_ (.A1(_06094_),
    .A2(_06343_),
    .B1(_05873_),
    .B2(_06344_),
    .C1(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__nand2_2 _20660_ (.A(_06345_),
    .B(_06347_),
    .Y(_06348_));
 sky130_vsdinv _20661_ (.A(_06348_),
    .Y(_06349_));
 sky130_vsdinv _20662_ (.A(_06342_),
    .Y(_06350_));
 sky130_fd_sc_hd__o22a_2 _20663_ (.A1(_06342_),
    .A2(_06349_),
    .B1(_06350_),
    .B2(_06348_),
    .X(_02643_));
 sky130_fd_sc_hd__o22a_2 _20664_ (.A1(_06336_),
    .A2(_06337_),
    .B1(_06099_),
    .B2(_06338_),
    .X(_06351_));
 sky130_fd_sc_hd__o22a_2 _20665_ (.A1(_06224_),
    .A2(_06268_),
    .B1(_06223_),
    .B2(_06269_),
    .X(_06352_));
 sky130_fd_sc_hd__o22a_2 _20666_ (.A1(_06246_),
    .A2(_06247_),
    .B1(_06225_),
    .B2(_06248_),
    .X(_06353_));
 sky130_fd_sc_hd__or2_2 _20667_ (.A(_06352_),
    .B(_06353_),
    .X(_06354_));
 sky130_fd_sc_hd__a21bo_2 _20668_ (.A1(_06352_),
    .A2(_06353_),
    .B1_N(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__o22a_2 _20669_ (.A1(_06265_),
    .A2(_06266_),
    .B1(_06249_),
    .B2(_06267_),
    .X(_06356_));
 sky130_fd_sc_hd__o22a_2 _20670_ (.A1(_06165_),
    .A2(_06327_),
    .B1(_06297_),
    .B2(_06328_),
    .X(_06357_));
 sky130_fd_sc_hd__a21oi_2 _20671_ (.A1(_06229_),
    .A2(_06230_),
    .B1(_06228_),
    .Y(_06358_));
 sky130_fd_sc_hd__buf_1 _20672_ (.A(_06110_),
    .X(_06359_));
 sky130_fd_sc_hd__buf_1 _20673_ (.A(_06359_),
    .X(_06360_));
 sky130_fd_sc_hd__buf_1 _20674_ (.A(_06232_),
    .X(_06361_));
 sky130_fd_sc_hd__buf_1 _20675_ (.A(_06361_),
    .X(_06362_));
 sky130_fd_sc_hd__o22a_2 _20676_ (.A1(_05702_),
    .A2(_06360_),
    .B1(_04695_),
    .B2(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__and4_2 _20677_ (.A(_11638_),
    .B(_11897_),
    .C(_11644_),
    .D(_11895_),
    .X(_06364_));
 sky130_fd_sc_hd__nor2_2 _20678_ (.A(_06363_),
    .B(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__nor2_2 _20679_ (.A(_06107_),
    .B(_06103_),
    .Y(_06366_));
 sky130_fd_sc_hd__a2bb2o_2 _20680_ (.A1_N(_06365_),
    .A2_N(_06366_),
    .B1(_06365_),
    .B2(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__buf_1 _20681_ (.A(_05826_),
    .X(_06368_));
 sky130_fd_sc_hd__buf_1 _20682_ (.A(_05827_),
    .X(_06369_));
 sky130_fd_sc_hd__o22a_2 _20683_ (.A1(_06368_),
    .A2(_06237_),
    .B1(_06369_),
    .B2(_05987_),
    .X(_06370_));
 sky130_fd_sc_hd__buf_1 _20684_ (.A(\pcpi_mul.rs1[21] ),
    .X(_06371_));
 sky130_fd_sc_hd__buf_1 _20685_ (.A(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__and4_2 _20686_ (.A(_11629_),
    .B(_06240_),
    .C(_11633_),
    .D(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__nor2_2 _20687_ (.A(_06370_),
    .B(_06373_),
    .Y(_06374_));
 sky130_vsdinv _20688_ (.A(\pcpi_mul.rs1[25] ),
    .Y(_06375_));
 sky130_fd_sc_hd__buf_1 _20689_ (.A(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__buf_1 _20690_ (.A(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__buf_1 _20691_ (.A(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__nor2_2 _20692_ (.A(_04538_),
    .B(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__a2bb2o_2 _20693_ (.A1_N(_06374_),
    .A2_N(_06379_),
    .B1(_06374_),
    .B2(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__o21ba_2 _20694_ (.A1(_06235_),
    .A2(_06242_),
    .B1_N(_06241_),
    .X(_06381_));
 sky130_fd_sc_hd__a2bb2o_2 _20695_ (.A1_N(_06380_),
    .A2_N(_06381_),
    .B1(_06380_),
    .B2(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__a2bb2o_2 _20696_ (.A1_N(_06367_),
    .A2_N(_06382_),
    .B1(_06367_),
    .B2(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__o22a_2 _20697_ (.A1(_06243_),
    .A2(_06244_),
    .B1(_06231_),
    .B2(_06245_),
    .X(_06384_));
 sky130_fd_sc_hd__a2bb2o_2 _20698_ (.A1_N(_06383_),
    .A2_N(_06384_),
    .B1(_06383_),
    .B2(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__a2bb2o_2 _20699_ (.A1_N(_06358_),
    .A2_N(_06385_),
    .B1(_06358_),
    .B2(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__o22a_2 _20700_ (.A1(_06253_),
    .A2(_06261_),
    .B1(_06252_),
    .B2(_06262_),
    .X(_06387_));
 sky130_fd_sc_hd__o22a_2 _20701_ (.A1(_06311_),
    .A2(_06312_),
    .B1(_06304_),
    .B2(_06313_),
    .X(_06388_));
 sky130_fd_sc_hd__o21ba_2 _20702_ (.A1(_06256_),
    .A2(_06260_),
    .B1_N(_06259_),
    .X(_06389_));
 sky130_fd_sc_hd__o21ba_2 _20703_ (.A1(_06298_),
    .A2(_06303_),
    .B1_N(_06302_),
    .X(_06390_));
 sky130_fd_sc_hd__or2_2 _20704_ (.A(_05735_),
    .B(_05815_),
    .X(_06391_));
 sky130_fd_sc_hd__buf_1 _20705_ (.A(\pcpi_mul.rs1[17] ),
    .X(_06392_));
 sky130_fd_sc_hd__buf_1 _20706_ (.A(\pcpi_mul.rs1[18] ),
    .X(_06393_));
 sky130_fd_sc_hd__and4_2 _20707_ (.A(_05742_),
    .B(_06392_),
    .C(_05744_),
    .D(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__o22a_2 _20708_ (.A1(_05738_),
    .A2(_05509_),
    .B1(_05739_),
    .B2(_06254_),
    .X(_06395_));
 sky130_fd_sc_hd__or2_2 _20709_ (.A(_06394_),
    .B(_06395_),
    .X(_06396_));
 sky130_fd_sc_hd__a2bb2o_2 _20710_ (.A1_N(_06391_),
    .A2_N(_06396_),
    .B1(_06391_),
    .B2(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__a2bb2o_2 _20711_ (.A1_N(_06390_),
    .A2_N(_06397_),
    .B1(_06390_),
    .B2(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__a2bb2o_2 _20712_ (.A1_N(_06389_),
    .A2_N(_06398_),
    .B1(_06389_),
    .B2(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__a2bb2o_2 _20713_ (.A1_N(_06388_),
    .A2_N(_06399_),
    .B1(_06388_),
    .B2(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__a2bb2o_2 _20714_ (.A1_N(_06387_),
    .A2_N(_06400_),
    .B1(_06387_),
    .B2(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__o22a_2 _20715_ (.A1(_06251_),
    .A2(_06263_),
    .B1(_06250_),
    .B2(_06264_),
    .X(_06402_));
 sky130_fd_sc_hd__a2bb2o_2 _20716_ (.A1_N(_06401_),
    .A2_N(_06402_),
    .B1(_06401_),
    .B2(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__a2bb2o_2 _20717_ (.A1_N(_06386_),
    .A2_N(_06403_),
    .B1(_06386_),
    .B2(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__a2bb2o_2 _20718_ (.A1_N(_06357_),
    .A2_N(_06404_),
    .B1(_06357_),
    .B2(_06404_),
    .X(_06405_));
 sky130_fd_sc_hd__a2bb2o_2 _20719_ (.A1_N(_06356_),
    .A2_N(_06405_),
    .B1(_06356_),
    .B2(_06405_),
    .X(_06406_));
 sky130_fd_sc_hd__o22a_2 _20720_ (.A1(_06324_),
    .A2(_06325_),
    .B1(_06314_),
    .B2(_06326_),
    .X(_06407_));
 sky130_fd_sc_hd__or2_2 _20721_ (.A(_06168_),
    .B(_05828_),
    .X(_06408_));
 sky130_fd_sc_hd__and4_2 _20722_ (.A(_06171_),
    .B(_05612_),
    .C(_06172_),
    .D(_06016_),
    .X(_06409_));
 sky130_fd_sc_hd__o22a_2 _20723_ (.A1(_05779_),
    .A2(_05255_),
    .B1(_06300_),
    .B2(_06014_),
    .X(_06410_));
 sky130_fd_sc_hd__or2_2 _20724_ (.A(_06409_),
    .B(_06410_),
    .X(_06411_));
 sky130_fd_sc_hd__a2bb2o_2 _20725_ (.A1_N(_06408_),
    .A2_N(_06411_),
    .B1(_06408_),
    .B2(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__or2_2 _20726_ (.A(_06176_),
    .B(_05736_),
    .X(_06413_));
 sky130_fd_sc_hd__and4_2 _20727_ (.A(_06182_),
    .B(_05433_),
    .C(_06183_),
    .D(_11924_),
    .X(_06414_));
 sky130_fd_sc_hd__buf_1 _20728_ (.A(_05130_),
    .X(_06415_));
 sky130_fd_sc_hd__o22a_2 _20729_ (.A1(_06307_),
    .A2(_05345_),
    .B1(_06415_),
    .B2(_05431_),
    .X(_06416_));
 sky130_fd_sc_hd__or2_2 _20730_ (.A(_06414_),
    .B(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__a2bb2o_2 _20731_ (.A1_N(_06413_),
    .A2_N(_06417_),
    .B1(_06413_),
    .B2(_06417_),
    .X(_06418_));
 sky130_fd_sc_hd__o21ba_2 _20732_ (.A1(_06306_),
    .A2(_06310_),
    .B1_N(_06309_),
    .X(_06419_));
 sky130_fd_sc_hd__a2bb2o_2 _20733_ (.A1_N(_06418_),
    .A2_N(_06419_),
    .B1(_06418_),
    .B2(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__a2bb2o_2 _20734_ (.A1_N(_06412_),
    .A2_N(_06420_),
    .B1(_06412_),
    .B2(_06420_),
    .X(_06421_));
 sky130_fd_sc_hd__o21ba_2 _20735_ (.A1(_06317_),
    .A2(_06321_),
    .B1_N(_06320_),
    .X(_06422_));
 sky130_fd_sc_hd__o21ba_2 _20736_ (.A1(_06278_),
    .A2(_06282_),
    .B1_N(_06281_),
    .X(_06423_));
 sky130_fd_sc_hd__or2_2 _20737_ (.A(_05309_),
    .B(_05164_),
    .X(_06424_));
 sky130_fd_sc_hd__buf_1 _20738_ (.A(_11601_),
    .X(_06425_));
 sky130_fd_sc_hd__buf_1 _20739_ (.A(_11604_),
    .X(_06426_));
 sky130_fd_sc_hd__and4_2 _20740_ (.A(_06425_),
    .B(_11934_),
    .C(_06426_),
    .D(_11931_),
    .X(_06427_));
 sky130_fd_sc_hd__buf_1 _20741_ (.A(_05795_),
    .X(_06428_));
 sky130_fd_sc_hd__buf_1 _20742_ (.A(_05013_),
    .X(_06429_));
 sky130_fd_sc_hd__o22a_2 _20743_ (.A1(_06428_),
    .A2(_05273_),
    .B1(_05388_),
    .B2(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__or2_2 _20744_ (.A(_06427_),
    .B(_06430_),
    .X(_06431_));
 sky130_fd_sc_hd__a2bb2o_2 _20745_ (.A1_N(_06424_),
    .A2_N(_06431_),
    .B1(_06424_),
    .B2(_06431_),
    .X(_06432_));
 sky130_fd_sc_hd__a2bb2o_2 _20746_ (.A1_N(_06423_),
    .A2_N(_06432_),
    .B1(_06423_),
    .B2(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__a2bb2o_2 _20747_ (.A1_N(_06422_),
    .A2_N(_06433_),
    .B1(_06422_),
    .B2(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__o22a_2 _20748_ (.A1(_06316_),
    .A2(_06322_),
    .B1(_06315_),
    .B2(_06323_),
    .X(_06435_));
 sky130_fd_sc_hd__a2bb2o_2 _20749_ (.A1_N(_06434_),
    .A2_N(_06435_),
    .B1(_06434_),
    .B2(_06435_),
    .X(_06436_));
 sky130_fd_sc_hd__a2bb2o_2 _20750_ (.A1_N(_06421_),
    .A2_N(_06436_),
    .B1(_06421_),
    .B2(_06436_),
    .X(_06437_));
 sky130_fd_sc_hd__a2bb2o_2 _20751_ (.A1_N(_06293_),
    .A2_N(_06437_),
    .B1(_06293_),
    .B2(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__a2bb2o_2 _20752_ (.A1_N(_06407_),
    .A2_N(_06438_),
    .B1(_06407_),
    .B2(_06438_),
    .X(_06439_));
 sky130_vsdinv _20753_ (.A(\pcpi_mul.rs2[25] ),
    .Y(_06440_));
 sky130_fd_sc_hd__buf_1 _20754_ (.A(_06440_),
    .X(_06441_));
 sky130_fd_sc_hd__buf_1 _20755_ (.A(_06441_),
    .X(_06442_));
 sky130_fd_sc_hd__buf_1 _20756_ (.A(_06442_),
    .X(_06443_));
 sky130_fd_sc_hd__o22a_2 _20757_ (.A1(_06443_),
    .A2(_04545_),
    .B1(_06275_),
    .B2(_04690_),
    .X(_06444_));
 sky130_fd_sc_hd__buf_1 _20758_ (.A(_06441_),
    .X(_06445_));
 sky130_fd_sc_hd__buf_1 _20759_ (.A(_06445_),
    .X(_06446_));
 sky130_fd_sc_hd__buf_1 _20760_ (.A(_06272_),
    .X(_06447_));
 sky130_fd_sc_hd__or4_2 _20761_ (.A(_06446_),
    .B(_04543_),
    .C(_06447_),
    .D(_04689_),
    .X(_06448_));
 sky130_fd_sc_hd__or2b_2 _20762_ (.A(_06444_),
    .B_N(_06448_),
    .X(_06449_));
 sky130_fd_sc_hd__o22a_2 _20763_ (.A1(_06288_),
    .A2(_06289_),
    .B1(_06283_),
    .B2(_06290_),
    .X(_06450_));
 sky130_fd_sc_hd__buf_1 _20764_ (.A(_05560_),
    .X(_06451_));
 sky130_fd_sc_hd__or2_2 _20765_ (.A(_06451_),
    .B(_05191_),
    .X(_06452_));
 sky130_fd_sc_hd__buf_1 _20766_ (.A(_11592_),
    .X(_06453_));
 sky130_fd_sc_hd__and4_2 _20767_ (.A(_06453_),
    .B(_11943_),
    .C(_06280_),
    .D(_05198_),
    .X(_06454_));
 sky130_fd_sc_hd__o22a_2 _20768_ (.A1(_06039_),
    .A2(_05194_),
    .B1(_05658_),
    .B2(_05312_),
    .X(_06455_));
 sky130_fd_sc_hd__or2_2 _20769_ (.A(_06454_),
    .B(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__a2bb2o_2 _20770_ (.A1_N(_06452_),
    .A2_N(_06456_),
    .B1(_06452_),
    .B2(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__or2_2 _20771_ (.A(_05925_),
    .B(_05137_),
    .X(_06458_));
 sky130_fd_sc_hd__and4_2 _20772_ (.A(_11584_),
    .B(_05144_),
    .C(\pcpi_mul.rs2[22] ),
    .D(_11948_),
    .X(_06459_));
 sky130_fd_sc_hd__o22a_2 _20773_ (.A1(_06158_),
    .A2(_04700_),
    .B1(_06029_),
    .B2(_04722_),
    .X(_06460_));
 sky130_fd_sc_hd__or2_2 _20774_ (.A(_06459_),
    .B(_06460_),
    .X(_06461_));
 sky130_fd_sc_hd__a2bb2o_2 _20775_ (.A1_N(_06458_),
    .A2_N(_06461_),
    .B1(_06458_),
    .B2(_06461_),
    .X(_06462_));
 sky130_fd_sc_hd__o21ba_2 _20776_ (.A1(_06284_),
    .A2(_06287_),
    .B1_N(_06286_),
    .X(_06463_));
 sky130_fd_sc_hd__a2bb2o_2 _20777_ (.A1_N(_06462_),
    .A2_N(_06463_),
    .B1(_06462_),
    .B2(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__a2bb2o_2 _20778_ (.A1_N(_06457_),
    .A2_N(_06464_),
    .B1(_06457_),
    .B2(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__or2_2 _20779_ (.A(_06450_),
    .B(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__a21bo_2 _20780_ (.A1(_06450_),
    .A2(_06465_),
    .B1_N(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__or2_2 _20781_ (.A(_06449_),
    .B(_06467_),
    .X(_06468_));
 sky130_fd_sc_hd__a21bo_2 _20782_ (.A1(_06449_),
    .A2(_06467_),
    .B1_N(_06468_),
    .X(_06469_));
 sky130_fd_sc_hd__a2bb2o_2 _20783_ (.A1_N(_06295_),
    .A2_N(_06469_),
    .B1(_06295_),
    .B2(_06469_),
    .X(_06470_));
 sky130_fd_sc_hd__a2bb2o_2 _20784_ (.A1_N(_06439_),
    .A2_N(_06470_),
    .B1(_06439_),
    .B2(_06470_),
    .X(_06471_));
 sky130_fd_sc_hd__a2bb2o_2 _20785_ (.A1_N(_06330_),
    .A2_N(_06471_),
    .B1(_06330_),
    .B2(_06471_),
    .X(_06472_));
 sky130_fd_sc_hd__a2bb2o_2 _20786_ (.A1_N(_06406_),
    .A2_N(_06472_),
    .B1(_06406_),
    .B2(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__o22a_2 _20787_ (.A1(_06205_),
    .A2(_06331_),
    .B1(_06270_),
    .B2(_06332_),
    .X(_06474_));
 sky130_fd_sc_hd__a2bb2o_2 _20788_ (.A1_N(_06473_),
    .A2_N(_06474_),
    .B1(_06473_),
    .B2(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__a2bb2o_2 _20789_ (.A1_N(_06355_),
    .A2_N(_06475_),
    .B1(_06355_),
    .B2(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__o22a_2 _20790_ (.A1(_06333_),
    .A2(_06334_),
    .B1(_06222_),
    .B2(_06335_),
    .X(_06477_));
 sky130_fd_sc_hd__a2bb2o_2 _20791_ (.A1_N(_06476_),
    .A2_N(_06477_),
    .B1(_06476_),
    .B2(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__a2bb2o_2 _20792_ (.A1_N(_06221_),
    .A2_N(_06478_),
    .B1(_06221_),
    .B2(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__or2_2 _20793_ (.A(_06351_),
    .B(_06479_),
    .X(_06480_));
 sky130_fd_sc_hd__a21bo_2 _20794_ (.A1(_06351_),
    .A2(_06479_),
    .B1_N(_06480_),
    .X(_06481_));
 sky130_fd_sc_hd__o21ai_2 _20795_ (.A1(_06342_),
    .A2(_06349_),
    .B1(_06341_),
    .Y(_06482_));
 sky130_fd_sc_hd__a2bb2o_2 _20796_ (.A1_N(_06481_),
    .A2_N(_06482_),
    .B1(_06481_),
    .B2(_06482_),
    .X(_02644_));
 sky130_fd_sc_hd__o22a_2 _20797_ (.A1(_06357_),
    .A2(_06404_),
    .B1(_06356_),
    .B2(_06405_),
    .X(_06483_));
 sky130_fd_sc_hd__o22a_2 _20798_ (.A1(_06383_),
    .A2(_06384_),
    .B1(_06358_),
    .B2(_06385_),
    .X(_06484_));
 sky130_fd_sc_hd__or2_2 _20799_ (.A(_06483_),
    .B(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__a21bo_2 _20800_ (.A1(_06483_),
    .A2(_06484_),
    .B1_N(_06485_),
    .X(_06486_));
 sky130_fd_sc_hd__o22a_2 _20801_ (.A1(_06401_),
    .A2(_06402_),
    .B1(_06386_),
    .B2(_06403_),
    .X(_06487_));
 sky130_fd_sc_hd__o22a_2 _20802_ (.A1(_06293_),
    .A2(_06437_),
    .B1(_06407_),
    .B2(_06438_),
    .X(_06488_));
 sky130_fd_sc_hd__a21oi_2 _20803_ (.A1(_06365_),
    .A2(_06366_),
    .B1(_06364_),
    .Y(_06489_));
 sky130_fd_sc_hd__o22a_2 _20804_ (.A1(_05702_),
    .A2(_06362_),
    .B1(_04695_),
    .B2(_06378_),
    .X(_06490_));
 sky130_fd_sc_hd__and4_2 _20805_ (.A(_11638_),
    .B(_11895_),
    .C(_11644_),
    .D(_11893_),
    .X(_06491_));
 sky130_fd_sc_hd__nor2_2 _20806_ (.A(_06490_),
    .B(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__nor2_2 _20807_ (.A(_06107_),
    .B(_06226_),
    .Y(_06493_));
 sky130_fd_sc_hd__a2bb2o_2 _20808_ (.A1_N(_06492_),
    .A2_N(_06493_),
    .B1(_06492_),
    .B2(_06493_),
    .X(_06494_));
 sky130_vsdinv _20809_ (.A(\pcpi_mul.rs1[26] ),
    .Y(_06495_));
 sky130_fd_sc_hd__buf_1 _20810_ (.A(_06495_),
    .X(_06496_));
 sky130_fd_sc_hd__buf_1 _20811_ (.A(_06496_),
    .X(_06497_));
 sky130_fd_sc_hd__or2_2 _20812_ (.A(_05713_),
    .B(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__buf_1 _20813_ (.A(\pcpi_mul.rs1[22] ),
    .X(_06499_));
 sky130_fd_sc_hd__and4_2 _20814_ (.A(_06115_),
    .B(_06372_),
    .C(_06116_),
    .D(_06499_),
    .X(_06500_));
 sky130_fd_sc_hd__buf_1 _20815_ (.A(_05891_),
    .X(_06501_));
 sky130_fd_sc_hd__buf_1 _20816_ (.A(_05994_),
    .X(_06502_));
 sky130_fd_sc_hd__o22a_2 _20817_ (.A1(_05718_),
    .A2(_06501_),
    .B1(_05719_),
    .B2(_06502_),
    .X(_06503_));
 sky130_fd_sc_hd__or2_2 _20818_ (.A(_06500_),
    .B(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__a2bb2o_2 _20819_ (.A1_N(_06498_),
    .A2_N(_06504_),
    .B1(_06498_),
    .B2(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__a21oi_2 _20820_ (.A1(_06374_),
    .A2(_06379_),
    .B1(_06373_),
    .Y(_06506_));
 sky130_fd_sc_hd__a2bb2o_2 _20821_ (.A1_N(_06505_),
    .A2_N(_06506_),
    .B1(_06505_),
    .B2(_06506_),
    .X(_06507_));
 sky130_fd_sc_hd__a2bb2o_2 _20822_ (.A1_N(_06494_),
    .A2_N(_06507_),
    .B1(_06494_),
    .B2(_06507_),
    .X(_06508_));
 sky130_fd_sc_hd__o22a_2 _20823_ (.A1(_06380_),
    .A2(_06381_),
    .B1(_06367_),
    .B2(_06382_),
    .X(_06509_));
 sky130_fd_sc_hd__a2bb2o_2 _20824_ (.A1_N(_06508_),
    .A2_N(_06509_),
    .B1(_06508_),
    .B2(_06509_),
    .X(_06510_));
 sky130_fd_sc_hd__a2bb2o_2 _20825_ (.A1_N(_06489_),
    .A2_N(_06510_),
    .B1(_06489_),
    .B2(_06510_),
    .X(_06511_));
 sky130_fd_sc_hd__o22a_2 _20826_ (.A1(_06390_),
    .A2(_06397_),
    .B1(_06389_),
    .B2(_06398_),
    .X(_06512_));
 sky130_fd_sc_hd__o22a_2 _20827_ (.A1(_06418_),
    .A2(_06419_),
    .B1(_06412_),
    .B2(_06420_),
    .X(_06513_));
 sky130_fd_sc_hd__o21ba_2 _20828_ (.A1(_06391_),
    .A2(_06396_),
    .B1_N(_06394_),
    .X(_06514_));
 sky130_fd_sc_hd__o21ba_2 _20829_ (.A1(_06408_),
    .A2(_06411_),
    .B1_N(_06409_),
    .X(_06515_));
 sky130_fd_sc_hd__or2_2 _20830_ (.A(_05735_),
    .B(_06237_),
    .X(_06516_));
 sky130_fd_sc_hd__buf_1 _20831_ (.A(\pcpi_mul.rs1[19] ),
    .X(_06517_));
 sky130_fd_sc_hd__and4_2 _20832_ (.A(_05742_),
    .B(_11910_),
    .C(_05744_),
    .D(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__o22a_2 _20833_ (.A1(_05738_),
    .A2(_05606_),
    .B1(_05739_),
    .B2(_05715_),
    .X(_06519_));
 sky130_fd_sc_hd__or2_2 _20834_ (.A(_06518_),
    .B(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__a2bb2o_2 _20835_ (.A1_N(_06516_),
    .A2_N(_06520_),
    .B1(_06516_),
    .B2(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__a2bb2o_2 _20836_ (.A1_N(_06515_),
    .A2_N(_06521_),
    .B1(_06515_),
    .B2(_06521_),
    .X(_06522_));
 sky130_fd_sc_hd__a2bb2o_2 _20837_ (.A1_N(_06514_),
    .A2_N(_06522_),
    .B1(_06514_),
    .B2(_06522_),
    .X(_06523_));
 sky130_fd_sc_hd__a2bb2o_2 _20838_ (.A1_N(_06513_),
    .A2_N(_06523_),
    .B1(_06513_),
    .B2(_06523_),
    .X(_06524_));
 sky130_fd_sc_hd__a2bb2o_2 _20839_ (.A1_N(_06512_),
    .A2_N(_06524_),
    .B1(_06512_),
    .B2(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__o22a_2 _20840_ (.A1(_06388_),
    .A2(_06399_),
    .B1(_06387_),
    .B2(_06400_),
    .X(_06526_));
 sky130_fd_sc_hd__a2bb2o_2 _20841_ (.A1_N(_06525_),
    .A2_N(_06526_),
    .B1(_06525_),
    .B2(_06526_),
    .X(_06527_));
 sky130_fd_sc_hd__a2bb2o_2 _20842_ (.A1_N(_06511_),
    .A2_N(_06527_),
    .B1(_06511_),
    .B2(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__a2bb2o_2 _20843_ (.A1_N(_06488_),
    .A2_N(_06528_),
    .B1(_06488_),
    .B2(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__a2bb2o_2 _20844_ (.A1_N(_06487_),
    .A2_N(_06529_),
    .B1(_06487_),
    .B2(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__o22a_2 _20845_ (.A1(_06434_),
    .A2(_06435_),
    .B1(_06421_),
    .B2(_06436_),
    .X(_06531_));
 sky130_fd_sc_hd__or2_2 _20846_ (.A(_06049_),
    .B(_05510_),
    .X(_06532_));
 sky130_fd_sc_hd__and4_2 _20847_ (.A(_06054_),
    .B(_06016_),
    .C(_06055_),
    .D(_11914_),
    .X(_06533_));
 sky130_fd_sc_hd__o22a_2 _20848_ (.A1(_06299_),
    .A2(_05342_),
    .B1(_06052_),
    .B2(_05501_),
    .X(_06534_));
 sky130_fd_sc_hd__or2_2 _20849_ (.A(_06533_),
    .B(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__a2bb2o_2 _20850_ (.A1_N(_06532_),
    .A2_N(_06535_),
    .B1(_06532_),
    .B2(_06535_),
    .X(_06536_));
 sky130_fd_sc_hd__or2_2 _20851_ (.A(_06305_),
    .B(_05845_),
    .X(_06537_));
 sky130_fd_sc_hd__and4_2 _20852_ (.A(_06182_),
    .B(_05514_),
    .C(_06183_),
    .D(_11922_),
    .X(_06538_));
 sky130_fd_sc_hd__o22a_2 _20853_ (.A1(_06307_),
    .A2(_05081_),
    .B1(_06179_),
    .B2(_05609_),
    .X(_06539_));
 sky130_fd_sc_hd__or2_2 _20854_ (.A(_06538_),
    .B(_06539_),
    .X(_06540_));
 sky130_fd_sc_hd__a2bb2o_2 _20855_ (.A1_N(_06537_),
    .A2_N(_06540_),
    .B1(_06537_),
    .B2(_06540_),
    .X(_06541_));
 sky130_fd_sc_hd__o21ba_2 _20856_ (.A1(_06413_),
    .A2(_06417_),
    .B1_N(_06414_),
    .X(_06542_));
 sky130_fd_sc_hd__a2bb2o_2 _20857_ (.A1_N(_06541_),
    .A2_N(_06542_),
    .B1(_06541_),
    .B2(_06542_),
    .X(_06543_));
 sky130_fd_sc_hd__a2bb2o_2 _20858_ (.A1_N(_06536_),
    .A2_N(_06543_),
    .B1(_06536_),
    .B2(_06543_),
    .X(_06544_));
 sky130_fd_sc_hd__o21ba_2 _20859_ (.A1(_06424_),
    .A2(_06431_),
    .B1_N(_06427_),
    .X(_06545_));
 sky130_fd_sc_hd__o21ba_2 _20860_ (.A1(_06452_),
    .A2(_06456_),
    .B1_N(_06454_),
    .X(_06546_));
 sky130_fd_sc_hd__or2_2 _20861_ (.A(_05309_),
    .B(_05155_),
    .X(_06547_));
 sky130_fd_sc_hd__and4_2 _20862_ (.A(_06425_),
    .B(_11931_),
    .C(_06426_),
    .D(_11929_),
    .X(_06548_));
 sky130_fd_sc_hd__buf_1 _20863_ (.A(_05391_),
    .X(_06549_));
 sky130_fd_sc_hd__o22a_2 _20864_ (.A1(_06428_),
    .A2(_06429_),
    .B1(_06549_),
    .B2(_06180_),
    .X(_06550_));
 sky130_fd_sc_hd__or2_2 _20865_ (.A(_06548_),
    .B(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__a2bb2o_2 _20866_ (.A1_N(_06547_),
    .A2_N(_06551_),
    .B1(_06547_),
    .B2(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__a2bb2o_2 _20867_ (.A1_N(_06546_),
    .A2_N(_06552_),
    .B1(_06546_),
    .B2(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__a2bb2o_2 _20868_ (.A1_N(_06545_),
    .A2_N(_06553_),
    .B1(_06545_),
    .B2(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__o22a_2 _20869_ (.A1(_06423_),
    .A2(_06432_),
    .B1(_06422_),
    .B2(_06433_),
    .X(_06555_));
 sky130_fd_sc_hd__a2bb2o_2 _20870_ (.A1_N(_06554_),
    .A2_N(_06555_),
    .B1(_06554_),
    .B2(_06555_),
    .X(_06556_));
 sky130_fd_sc_hd__a2bb2o_2 _20871_ (.A1_N(_06544_),
    .A2_N(_06556_),
    .B1(_06544_),
    .B2(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__a2bb2o_2 _20872_ (.A1_N(_06466_),
    .A2_N(_06557_),
    .B1(_06466_),
    .B2(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__a2bb2o_2 _20873_ (.A1_N(_06531_),
    .A2_N(_06558_),
    .B1(_06531_),
    .B2(_06558_),
    .X(_06559_));
 sky130_fd_sc_hd__or2_2 _20874_ (.A(_06271_),
    .B(_05061_),
    .X(_06560_));
 sky130_fd_sc_hd__and4_2 _20875_ (.A(_11579_),
    .B(_11954_),
    .C(\pcpi_mul.rs2[26] ),
    .D(_11956_),
    .X(_06561_));
 sky130_vsdinv _20876_ (.A(\pcpi_mul.rs2[26] ),
    .Y(_06562_));
 sky130_fd_sc_hd__o22a_2 _20877_ (.A1(_06440_),
    .A2(_04687_),
    .B1(_06562_),
    .B2(_04541_),
    .X(_06563_));
 sky130_fd_sc_hd__or2_2 _20878_ (.A(_06561_),
    .B(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__a2bb2o_2 _20879_ (.A1_N(_06560_),
    .A2_N(_06564_),
    .B1(_06560_),
    .B2(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__or2_2 _20880_ (.A(_06448_),
    .B(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__a21bo_2 _20881_ (.A1(_06448_),
    .A2(_06565_),
    .B1_N(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__buf_1 _20882_ (.A(_05086_),
    .X(_06568_));
 sky130_fd_sc_hd__or2_2 _20883_ (.A(_06451_),
    .B(_06568_),
    .X(_06569_));
 sky130_fd_sc_hd__buf_1 _20884_ (.A(_11597_),
    .X(_06570_));
 sky130_fd_sc_hd__and4_2 _20885_ (.A(_06453_),
    .B(_11940_),
    .C(_06570_),
    .D(_05577_),
    .X(_06571_));
 sky130_fd_sc_hd__buf_1 _20886_ (.A(_05773_),
    .X(_06572_));
 sky130_fd_sc_hd__buf_1 _20887_ (.A(_05657_),
    .X(_06573_));
 sky130_fd_sc_hd__o22a_2 _20888_ (.A1(_06572_),
    .A2(_05195_),
    .B1(_06573_),
    .B2(_05396_),
    .X(_06574_));
 sky130_fd_sc_hd__or2_2 _20889_ (.A(_06571_),
    .B(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__a2bb2o_2 _20890_ (.A1_N(_06569_),
    .A2_N(_06575_),
    .B1(_06569_),
    .B2(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__or2_2 _20891_ (.A(_05925_),
    .B(_05225_),
    .X(_06577_));
 sky130_fd_sc_hd__and4_2 _20892_ (.A(_11584_),
    .B(_05145_),
    .C(_11588_),
    .D(_05316_),
    .X(_06578_));
 sky130_fd_sc_hd__buf_1 _20893_ (.A(_06158_),
    .X(_06579_));
 sky130_fd_sc_hd__o22a_2 _20894_ (.A1(_06579_),
    .A2(_04722_),
    .B1(_06029_),
    .B2(_04975_),
    .X(_06580_));
 sky130_fd_sc_hd__or2_2 _20895_ (.A(_06578_),
    .B(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__a2bb2o_2 _20896_ (.A1_N(_06577_),
    .A2_N(_06581_),
    .B1(_06577_),
    .B2(_06581_),
    .X(_06582_));
 sky130_fd_sc_hd__o21ba_2 _20897_ (.A1(_06458_),
    .A2(_06461_),
    .B1_N(_06459_),
    .X(_06583_));
 sky130_fd_sc_hd__a2bb2o_2 _20898_ (.A1_N(_06582_),
    .A2_N(_06583_),
    .B1(_06582_),
    .B2(_06583_),
    .X(_06584_));
 sky130_fd_sc_hd__a2bb2o_2 _20899_ (.A1_N(_06576_),
    .A2_N(_06584_),
    .B1(_06576_),
    .B2(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__o22a_2 _20900_ (.A1(_06462_),
    .A2(_06463_),
    .B1(_06457_),
    .B2(_06464_),
    .X(_06586_));
 sky130_fd_sc_hd__or2_2 _20901_ (.A(_06585_),
    .B(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__a21bo_2 _20902_ (.A1(_06585_),
    .A2(_06586_),
    .B1_N(_06587_),
    .X(_06588_));
 sky130_fd_sc_hd__or2_2 _20903_ (.A(_06567_),
    .B(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__a21bo_2 _20904_ (.A1(_06567_),
    .A2(_06588_),
    .B1_N(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__a2bb2o_2 _20905_ (.A1_N(_06468_),
    .A2_N(_06590_),
    .B1(_06468_),
    .B2(_06590_),
    .X(_06591_));
 sky130_fd_sc_hd__a2bb2o_2 _20906_ (.A1_N(_06559_),
    .A2_N(_06591_),
    .B1(_06559_),
    .B2(_06591_),
    .X(_06592_));
 sky130_fd_sc_hd__o22a_2 _20907_ (.A1(_06295_),
    .A2(_06469_),
    .B1(_06439_),
    .B2(_06470_),
    .X(_06593_));
 sky130_fd_sc_hd__a2bb2o_2 _20908_ (.A1_N(_06592_),
    .A2_N(_06593_),
    .B1(_06592_),
    .B2(_06593_),
    .X(_06594_));
 sky130_fd_sc_hd__a2bb2o_2 _20909_ (.A1_N(_06530_),
    .A2_N(_06594_),
    .B1(_06530_),
    .B2(_06594_),
    .X(_06595_));
 sky130_fd_sc_hd__o22a_2 _20910_ (.A1(_06330_),
    .A2(_06471_),
    .B1(_06406_),
    .B2(_06472_),
    .X(_06596_));
 sky130_fd_sc_hd__a2bb2o_2 _20911_ (.A1_N(_06595_),
    .A2_N(_06596_),
    .B1(_06595_),
    .B2(_06596_),
    .X(_06597_));
 sky130_fd_sc_hd__a2bb2o_2 _20912_ (.A1_N(_06486_),
    .A2_N(_06597_),
    .B1(_06486_),
    .B2(_06597_),
    .X(_06598_));
 sky130_fd_sc_hd__o22a_2 _20913_ (.A1(_06473_),
    .A2(_06474_),
    .B1(_06355_),
    .B2(_06475_),
    .X(_06599_));
 sky130_fd_sc_hd__a2bb2o_2 _20914_ (.A1_N(_06598_),
    .A2_N(_06599_),
    .B1(_06598_),
    .B2(_06599_),
    .X(_06600_));
 sky130_fd_sc_hd__a2bb2o_2 _20915_ (.A1_N(_06354_),
    .A2_N(_06600_),
    .B1(_06354_),
    .B2(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__o22a_2 _20916_ (.A1(_06476_),
    .A2(_06477_),
    .B1(_06221_),
    .B2(_06478_),
    .X(_06602_));
 sky130_fd_sc_hd__or2_2 _20917_ (.A(_06601_),
    .B(_06602_),
    .X(_06603_));
 sky130_fd_sc_hd__a21bo_2 _20918_ (.A1(_06601_),
    .A2(_06602_),
    .B1_N(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__a22o_2 _20919_ (.A1(_06351_),
    .A2(_06479_),
    .B1(_06341_),
    .B2(_06480_),
    .X(_06605_));
 sky130_fd_sc_hd__o31a_2 _20920_ (.A1(_06342_),
    .A2(_06481_),
    .A3(_06349_),
    .B1(_06605_),
    .X(_06606_));
 sky130_fd_sc_hd__a2bb2oi_2 _20921_ (.A1_N(_06604_),
    .A2_N(_06606_),
    .B1(_06604_),
    .B2(_06606_),
    .Y(_02645_));
 sky130_fd_sc_hd__o22a_2 _20922_ (.A1(_06598_),
    .A2(_06599_),
    .B1(_06354_),
    .B2(_06600_),
    .X(_06607_));
 sky130_fd_sc_hd__o22a_2 _20923_ (.A1(_06488_),
    .A2(_06528_),
    .B1(_06487_),
    .B2(_06529_),
    .X(_06608_));
 sky130_fd_sc_hd__o22a_2 _20924_ (.A1(_06508_),
    .A2(_06509_),
    .B1(_06489_),
    .B2(_06510_),
    .X(_06609_));
 sky130_fd_sc_hd__or2_2 _20925_ (.A(_06608_),
    .B(_06609_),
    .X(_06610_));
 sky130_fd_sc_hd__a21bo_2 _20926_ (.A1(_06608_),
    .A2(_06609_),
    .B1_N(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__o22a_2 _20927_ (.A1(_06525_),
    .A2(_06526_),
    .B1(_06511_),
    .B2(_06527_),
    .X(_06612_));
 sky130_fd_sc_hd__o22a_2 _20928_ (.A1(_06466_),
    .A2(_06557_),
    .B1(_06531_),
    .B2(_06558_),
    .X(_06613_));
 sky130_fd_sc_hd__a21oi_2 _20929_ (.A1(_06492_),
    .A2(_06493_),
    .B1(_06491_),
    .Y(_06614_));
 sky130_fd_sc_hd__and4_2 _20930_ (.A(_11637_),
    .B(_11893_),
    .C(_11643_),
    .D(_11889_),
    .X(_06615_));
 sky130_fd_sc_hd__buf_1 _20931_ (.A(_06375_),
    .X(_06616_));
 sky130_fd_sc_hd__buf_1 _20932_ (.A(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__o22a_2 _20933_ (.A1(_05813_),
    .A2(_06617_),
    .B1(_05156_),
    .B2(_06497_),
    .X(_06618_));
 sky130_fd_sc_hd__or2_2 _20934_ (.A(_06615_),
    .B(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__buf_1 _20935_ (.A(_06234_),
    .X(_06620_));
 sky130_fd_sc_hd__or2_2 _20936_ (.A(_05162_),
    .B(_06620_),
    .X(_06621_));
 sky130_fd_sc_hd__a2bb2o_2 _20937_ (.A1_N(_06619_),
    .A2_N(_06621_),
    .B1(_06619_),
    .B2(_06621_),
    .X(_06622_));
 sky130_vsdinv _20938_ (.A(\pcpi_mul.rs1[27] ),
    .Y(_06623_));
 sky130_fd_sc_hd__buf_1 _20939_ (.A(_06623_),
    .X(_06624_));
 sky130_fd_sc_hd__buf_1 _20940_ (.A(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__or2_2 _20941_ (.A(_05713_),
    .B(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__buf_1 _20942_ (.A(\pcpi_mul.rs1[23] ),
    .X(_06627_));
 sky130_fd_sc_hd__and4_2 _20943_ (.A(_06115_),
    .B(_11900_),
    .C(_06116_),
    .D(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__o22a_2 _20944_ (.A1(_05718_),
    .A2(_06502_),
    .B1(_05719_),
    .B2(_06359_),
    .X(_06629_));
 sky130_fd_sc_hd__or2_2 _20945_ (.A(_06628_),
    .B(_06629_),
    .X(_06630_));
 sky130_fd_sc_hd__a2bb2o_2 _20946_ (.A1_N(_06626_),
    .A2_N(_06630_),
    .B1(_06626_),
    .B2(_06630_),
    .X(_06631_));
 sky130_fd_sc_hd__o21ba_2 _20947_ (.A1(_06498_),
    .A2(_06504_),
    .B1_N(_06500_),
    .X(_06632_));
 sky130_fd_sc_hd__a2bb2o_2 _20948_ (.A1_N(_06631_),
    .A2_N(_06632_),
    .B1(_06631_),
    .B2(_06632_),
    .X(_06633_));
 sky130_fd_sc_hd__a2bb2o_2 _20949_ (.A1_N(_06622_),
    .A2_N(_06633_),
    .B1(_06622_),
    .B2(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__o22a_2 _20950_ (.A1(_06505_),
    .A2(_06506_),
    .B1(_06494_),
    .B2(_06507_),
    .X(_06635_));
 sky130_fd_sc_hd__a2bb2o_2 _20951_ (.A1_N(_06634_),
    .A2_N(_06635_),
    .B1(_06634_),
    .B2(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__a2bb2o_2 _20952_ (.A1_N(_06614_),
    .A2_N(_06636_),
    .B1(_06614_),
    .B2(_06636_),
    .X(_06637_));
 sky130_fd_sc_hd__o22a_2 _20953_ (.A1(_06515_),
    .A2(_06521_),
    .B1(_06514_),
    .B2(_06522_),
    .X(_06638_));
 sky130_fd_sc_hd__o22a_2 _20954_ (.A1(_06541_),
    .A2(_06542_),
    .B1(_06536_),
    .B2(_06543_),
    .X(_06639_));
 sky130_fd_sc_hd__o21ba_2 _20955_ (.A1(_06516_),
    .A2(_06520_),
    .B1_N(_06518_),
    .X(_06640_));
 sky130_fd_sc_hd__o21ba_2 _20956_ (.A1(_06532_),
    .A2(_06535_),
    .B1_N(_06533_),
    .X(_06641_));
 sky130_fd_sc_hd__or2_2 _20957_ (.A(_05735_),
    .B(_05987_),
    .X(_06642_));
 sky130_fd_sc_hd__and4_2 _20958_ (.A(_06136_),
    .B(_11908_),
    .C(_06137_),
    .D(_06239_),
    .X(_06643_));
 sky130_fd_sc_hd__o22a_2 _20959_ (.A1(_05738_),
    .A2(_05814_),
    .B1(_05739_),
    .B2(_06236_),
    .X(_06644_));
 sky130_fd_sc_hd__or2_2 _20960_ (.A(_06643_),
    .B(_06644_),
    .X(_06645_));
 sky130_fd_sc_hd__a2bb2o_2 _20961_ (.A1_N(_06642_),
    .A2_N(_06645_),
    .B1(_06642_),
    .B2(_06645_),
    .X(_06646_));
 sky130_fd_sc_hd__a2bb2o_2 _20962_ (.A1_N(_06641_),
    .A2_N(_06646_),
    .B1(_06641_),
    .B2(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__a2bb2o_2 _20963_ (.A1_N(_06640_),
    .A2_N(_06647_),
    .B1(_06640_),
    .B2(_06647_),
    .X(_06648_));
 sky130_fd_sc_hd__a2bb2o_2 _20964_ (.A1_N(_06639_),
    .A2_N(_06648_),
    .B1(_06639_),
    .B2(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__a2bb2o_2 _20965_ (.A1_N(_06638_),
    .A2_N(_06649_),
    .B1(_06638_),
    .B2(_06649_),
    .X(_06650_));
 sky130_fd_sc_hd__o22a_2 _20966_ (.A1(_06513_),
    .A2(_06523_),
    .B1(_06512_),
    .B2(_06524_),
    .X(_06651_));
 sky130_fd_sc_hd__a2bb2o_2 _20967_ (.A1_N(_06650_),
    .A2_N(_06651_),
    .B1(_06650_),
    .B2(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__a2bb2o_2 _20968_ (.A1_N(_06637_),
    .A2_N(_06652_),
    .B1(_06637_),
    .B2(_06652_),
    .X(_06653_));
 sky130_fd_sc_hd__a2bb2o_2 _20969_ (.A1_N(_06613_),
    .A2_N(_06653_),
    .B1(_06613_),
    .B2(_06653_),
    .X(_06654_));
 sky130_fd_sc_hd__a2bb2o_2 _20970_ (.A1_N(_06612_),
    .A2_N(_06654_),
    .B1(_06612_),
    .B2(_06654_),
    .X(_06655_));
 sky130_fd_sc_hd__o22a_2 _20971_ (.A1(_06554_),
    .A2(_06555_),
    .B1(_06544_),
    .B2(_06556_),
    .X(_06656_));
 sky130_fd_sc_hd__or2_2 _20972_ (.A(_06168_),
    .B(_06255_),
    .X(_06657_));
 sky130_fd_sc_hd__and4_2 _20973_ (.A(_06054_),
    .B(_11914_),
    .C(_06055_),
    .D(_11912_),
    .X(_06658_));
 sky130_fd_sc_hd__o22a_2 _20974_ (.A1(_06299_),
    .A2(_05428_),
    .B1(_06300_),
    .B2(_06257_),
    .X(_06659_));
 sky130_fd_sc_hd__or2_2 _20975_ (.A(_06658_),
    .B(_06659_),
    .X(_06660_));
 sky130_fd_sc_hd__a2bb2o_2 _20976_ (.A1_N(_06657_),
    .A2_N(_06660_),
    .B1(_06657_),
    .B2(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__or2_2 _20977_ (.A(_06305_),
    .B(_05720_),
    .X(_06662_));
 sky130_fd_sc_hd__and4_2 _20978_ (.A(_06182_),
    .B(_11922_),
    .C(_06183_),
    .D(_05612_),
    .X(_06663_));
 sky130_fd_sc_hd__o22a_2 _20979_ (.A1(_06307_),
    .A2(_05168_),
    .B1(_06179_),
    .B2(_05610_),
    .X(_06664_));
 sky130_fd_sc_hd__or2_2 _20980_ (.A(_06663_),
    .B(_06664_),
    .X(_06665_));
 sky130_fd_sc_hd__a2bb2o_2 _20981_ (.A1_N(_06662_),
    .A2_N(_06665_),
    .B1(_06662_),
    .B2(_06665_),
    .X(_06666_));
 sky130_fd_sc_hd__o21ba_2 _20982_ (.A1(_06537_),
    .A2(_06540_),
    .B1_N(_06538_),
    .X(_06667_));
 sky130_fd_sc_hd__a2bb2o_2 _20983_ (.A1_N(_06666_),
    .A2_N(_06667_),
    .B1(_06666_),
    .B2(_06667_),
    .X(_06668_));
 sky130_fd_sc_hd__a2bb2o_2 _20984_ (.A1_N(_06661_),
    .A2_N(_06668_),
    .B1(_06661_),
    .B2(_06668_),
    .X(_06669_));
 sky130_fd_sc_hd__o21ba_2 _20985_ (.A1(_06547_),
    .A2(_06551_),
    .B1_N(_06548_),
    .X(_06670_));
 sky130_fd_sc_hd__o21ba_2 _20986_ (.A1(_06569_),
    .A2(_06575_),
    .B1_N(_06571_),
    .X(_06671_));
 sky130_fd_sc_hd__or2_2 _20987_ (.A(_05309_),
    .B(_05937_),
    .X(_06672_));
 sky130_fd_sc_hd__and4_2 _20988_ (.A(_06425_),
    .B(_06184_),
    .C(_06426_),
    .D(_05743_),
    .X(_06673_));
 sky130_fd_sc_hd__o22a_2 _20989_ (.A1(_06428_),
    .A2(_05258_),
    .B1(_06549_),
    .B2(_05530_),
    .X(_06674_));
 sky130_fd_sc_hd__or2_2 _20990_ (.A(_06673_),
    .B(_06674_),
    .X(_06675_));
 sky130_fd_sc_hd__a2bb2o_2 _20991_ (.A1_N(_06672_),
    .A2_N(_06675_),
    .B1(_06672_),
    .B2(_06675_),
    .X(_06676_));
 sky130_fd_sc_hd__a2bb2o_2 _20992_ (.A1_N(_06671_),
    .A2_N(_06676_),
    .B1(_06671_),
    .B2(_06676_),
    .X(_06677_));
 sky130_fd_sc_hd__a2bb2o_2 _20993_ (.A1_N(_06670_),
    .A2_N(_06677_),
    .B1(_06670_),
    .B2(_06677_),
    .X(_06678_));
 sky130_fd_sc_hd__o22a_2 _20994_ (.A1(_06546_),
    .A2(_06552_),
    .B1(_06545_),
    .B2(_06553_),
    .X(_06679_));
 sky130_fd_sc_hd__a2bb2o_2 _20995_ (.A1_N(_06678_),
    .A2_N(_06679_),
    .B1(_06678_),
    .B2(_06679_),
    .X(_06680_));
 sky130_fd_sc_hd__a2bb2o_2 _20996_ (.A1_N(_06669_),
    .A2_N(_06680_),
    .B1(_06669_),
    .B2(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__a2bb2o_2 _20997_ (.A1_N(_06587_),
    .A2_N(_06681_),
    .B1(_06587_),
    .B2(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__a2bb2o_2 _20998_ (.A1_N(_06656_),
    .A2_N(_06682_),
    .B1(_06656_),
    .B2(_06682_),
    .X(_06683_));
 sky130_vsdinv _20999_ (.A(\pcpi_mul.rs2[27] ),
    .Y(_06684_));
 sky130_fd_sc_hd__buf_1 _21000_ (.A(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__buf_1 _21001_ (.A(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__buf_1 _21002_ (.A(_06686_),
    .X(_06687_));
 sky130_fd_sc_hd__or2_2 _21003_ (.A(_06687_),
    .B(_04544_),
    .X(_06688_));
 sky130_fd_sc_hd__or2_2 _21004_ (.A(_06271_),
    .B(_05406_),
    .X(_06689_));
 sky130_fd_sc_hd__o22a_2 _21005_ (.A1(_06562_),
    .A2(_04751_),
    .B1(_06440_),
    .B2(_04701_),
    .X(_06690_));
 sky130_fd_sc_hd__and4_2 _21006_ (.A(\pcpi_mul.rs2[26] ),
    .B(_05238_),
    .C(\pcpi_mul.rs2[25] ),
    .D(_11951_),
    .X(_06691_));
 sky130_fd_sc_hd__or2_2 _21007_ (.A(_06690_),
    .B(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__a2bb2o_2 _21008_ (.A1_N(_06689_),
    .A2_N(_06692_),
    .B1(_06689_),
    .B2(_06692_),
    .X(_06693_));
 sky130_fd_sc_hd__o21ba_2 _21009_ (.A1(_06560_),
    .A2(_06564_),
    .B1_N(_06561_),
    .X(_06694_));
 sky130_fd_sc_hd__or2_2 _21010_ (.A(_06693_),
    .B(_06694_),
    .X(_06695_));
 sky130_fd_sc_hd__a21bo_2 _21011_ (.A1(_06693_),
    .A2(_06694_),
    .B1_N(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__or2_2 _21012_ (.A(_06688_),
    .B(_06696_),
    .X(_06697_));
 sky130_fd_sc_hd__a21bo_2 _21013_ (.A1(_06688_),
    .A2(_06696_),
    .B1_N(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__o22a_2 _21014_ (.A1(_06582_),
    .A2(_06583_),
    .B1(_06576_),
    .B2(_06584_),
    .X(_06699_));
 sky130_fd_sc_hd__buf_1 _21015_ (.A(_05561_),
    .X(_06700_));
 sky130_fd_sc_hd__or2_2 _21016_ (.A(_06700_),
    .B(_05077_),
    .X(_06701_));
 sky130_fd_sc_hd__o22a_2 _21017_ (.A1(_06572_),
    .A2(_05575_),
    .B1(_06573_),
    .B2(_05273_),
    .X(_06702_));
 sky130_fd_sc_hd__buf_1 _21018_ (.A(_11592_),
    .X(_06703_));
 sky130_fd_sc_hd__and4_2 _21019_ (.A(_06703_),
    .B(_11937_),
    .C(_06570_),
    .D(_05176_),
    .X(_06704_));
 sky130_fd_sc_hd__or2_2 _21020_ (.A(_06702_),
    .B(_06704_),
    .X(_06705_));
 sky130_fd_sc_hd__a2bb2o_2 _21021_ (.A1_N(_06701_),
    .A2_N(_06705_),
    .B1(_06701_),
    .B2(_06705_),
    .X(_06706_));
 sky130_fd_sc_hd__or2_2 _21022_ (.A(_06035_),
    .B(_05312_),
    .X(_06707_));
 sky130_fd_sc_hd__and4_2 _21023_ (.A(_11584_),
    .B(_05316_),
    .C(_11588_),
    .D(_05197_),
    .X(_06708_));
 sky130_fd_sc_hd__o22a_2 _21024_ (.A1(_06579_),
    .A2(_05227_),
    .B1(_06033_),
    .B2(_05194_),
    .X(_06709_));
 sky130_fd_sc_hd__or2_2 _21025_ (.A(_06708_),
    .B(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__a2bb2o_2 _21026_ (.A1_N(_06707_),
    .A2_N(_06710_),
    .B1(_06707_),
    .B2(_06710_),
    .X(_06711_));
 sky130_fd_sc_hd__o21ba_2 _21027_ (.A1(_06577_),
    .A2(_06581_),
    .B1_N(_06578_),
    .X(_06712_));
 sky130_fd_sc_hd__a2bb2o_2 _21028_ (.A1_N(_06711_),
    .A2_N(_06712_),
    .B1(_06711_),
    .B2(_06712_),
    .X(_06713_));
 sky130_fd_sc_hd__a2bb2o_2 _21029_ (.A1_N(_06706_),
    .A2_N(_06713_),
    .B1(_06706_),
    .B2(_06713_),
    .X(_06714_));
 sky130_fd_sc_hd__a2bb2o_2 _21030_ (.A1_N(_06566_),
    .A2_N(_06714_),
    .B1(_06566_),
    .B2(_06714_),
    .X(_06715_));
 sky130_fd_sc_hd__a2bb2o_2 _21031_ (.A1_N(_06699_),
    .A2_N(_06715_),
    .B1(_06699_),
    .B2(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__or2_2 _21032_ (.A(_06698_),
    .B(_06716_),
    .X(_06717_));
 sky130_fd_sc_hd__a21bo_2 _21033_ (.A1(_06698_),
    .A2(_06716_),
    .B1_N(_06717_),
    .X(_06718_));
 sky130_fd_sc_hd__a2bb2o_2 _21034_ (.A1_N(_06589_),
    .A2_N(_06718_),
    .B1(_06589_),
    .B2(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__a2bb2o_2 _21035_ (.A1_N(_06683_),
    .A2_N(_06719_),
    .B1(_06683_),
    .B2(_06719_),
    .X(_06720_));
 sky130_fd_sc_hd__o22a_2 _21036_ (.A1(_06468_),
    .A2(_06590_),
    .B1(_06559_),
    .B2(_06591_),
    .X(_06721_));
 sky130_fd_sc_hd__a2bb2o_2 _21037_ (.A1_N(_06720_),
    .A2_N(_06721_),
    .B1(_06720_),
    .B2(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__a2bb2o_2 _21038_ (.A1_N(_06655_),
    .A2_N(_06722_),
    .B1(_06655_),
    .B2(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__o22a_2 _21039_ (.A1(_06592_),
    .A2(_06593_),
    .B1(_06530_),
    .B2(_06594_),
    .X(_06724_));
 sky130_fd_sc_hd__a2bb2o_2 _21040_ (.A1_N(_06723_),
    .A2_N(_06724_),
    .B1(_06723_),
    .B2(_06724_),
    .X(_06725_));
 sky130_fd_sc_hd__a2bb2o_2 _21041_ (.A1_N(_06611_),
    .A2_N(_06725_),
    .B1(_06611_),
    .B2(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__o22a_2 _21042_ (.A1(_06595_),
    .A2(_06596_),
    .B1(_06486_),
    .B2(_06597_),
    .X(_06727_));
 sky130_fd_sc_hd__a2bb2o_2 _21043_ (.A1_N(_06726_),
    .A2_N(_06727_),
    .B1(_06726_),
    .B2(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__a2bb2o_2 _21044_ (.A1_N(_06485_),
    .A2_N(_06728_),
    .B1(_06485_),
    .B2(_06728_),
    .X(_06729_));
 sky130_fd_sc_hd__and2_2 _21045_ (.A(_06607_),
    .B(_06729_),
    .X(_06730_));
 sky130_fd_sc_hd__or2_2 _21046_ (.A(_06607_),
    .B(_06729_),
    .X(_06731_));
 sky130_fd_sc_hd__or2b_2 _21047_ (.A(_06730_),
    .B_N(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__o21ai_2 _21048_ (.A1(_06604_),
    .A2(_06606_),
    .B1(_06603_),
    .Y(_06733_));
 sky130_fd_sc_hd__a2bb2o_2 _21049_ (.A1_N(_06732_),
    .A2_N(_06733_),
    .B1(_06732_),
    .B2(_06733_),
    .X(_02646_));
 sky130_fd_sc_hd__o22a_2 _21050_ (.A1(_06613_),
    .A2(_06653_),
    .B1(_06612_),
    .B2(_06654_),
    .X(_06734_));
 sky130_fd_sc_hd__o22a_2 _21051_ (.A1(_06634_),
    .A2(_06635_),
    .B1(_06614_),
    .B2(_06636_),
    .X(_06735_));
 sky130_fd_sc_hd__or2_2 _21052_ (.A(_06734_),
    .B(_06735_),
    .X(_06736_));
 sky130_fd_sc_hd__a21bo_2 _21053_ (.A1(_06734_),
    .A2(_06735_),
    .B1_N(_06736_),
    .X(_06737_));
 sky130_fd_sc_hd__o22a_2 _21054_ (.A1(_06650_),
    .A2(_06651_),
    .B1(_06637_),
    .B2(_06652_),
    .X(_06738_));
 sky130_fd_sc_hd__o22a_2 _21055_ (.A1(_06587_),
    .A2(_06681_),
    .B1(_06656_),
    .B2(_06682_),
    .X(_06739_));
 sky130_fd_sc_hd__o21ba_2 _21056_ (.A1(_06619_),
    .A2(_06621_),
    .B1_N(_06615_),
    .X(_06740_));
 sky130_fd_sc_hd__and4_2 _21057_ (.A(_11637_),
    .B(_11889_),
    .C(_11643_),
    .D(_11885_),
    .X(_06741_));
 sky130_fd_sc_hd__buf_1 _21058_ (.A(_06495_),
    .X(_06742_));
 sky130_fd_sc_hd__buf_1 _21059_ (.A(_06742_),
    .X(_06743_));
 sky130_fd_sc_hd__o22a_2 _21060_ (.A1(_05153_),
    .A2(_06743_),
    .B1(_05156_),
    .B2(_06625_),
    .X(_06744_));
 sky130_fd_sc_hd__or2_2 _21061_ (.A(_06741_),
    .B(_06744_),
    .X(_06745_));
 sky130_fd_sc_hd__or2_2 _21062_ (.A(_05162_),
    .B(_06378_),
    .X(_06746_));
 sky130_fd_sc_hd__a2bb2o_2 _21063_ (.A1_N(_06745_),
    .A2_N(_06746_),
    .B1(_06745_),
    .B2(_06746_),
    .X(_06747_));
 sky130_vsdinv _21064_ (.A(\pcpi_mul.rs1[28] ),
    .Y(_06748_));
 sky130_fd_sc_hd__buf_1 _21065_ (.A(_06748_),
    .X(_06749_));
 sky130_fd_sc_hd__buf_1 _21066_ (.A(_06749_),
    .X(_06750_));
 sky130_fd_sc_hd__or2_2 _21067_ (.A(_05713_),
    .B(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__buf_1 _21068_ (.A(\pcpi_mul.rs1[24] ),
    .X(_06752_));
 sky130_fd_sc_hd__and4_2 _21069_ (.A(_06115_),
    .B(_06627_),
    .C(_06116_),
    .D(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__buf_1 _21070_ (.A(_06110_),
    .X(_06754_));
 sky130_fd_sc_hd__o22a_2 _21071_ (.A1(_05718_),
    .A2(_06754_),
    .B1(_05719_),
    .B2(_06361_),
    .X(_06755_));
 sky130_fd_sc_hd__or2_2 _21072_ (.A(_06753_),
    .B(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__a2bb2o_2 _21073_ (.A1_N(_06751_),
    .A2_N(_06756_),
    .B1(_06751_),
    .B2(_06756_),
    .X(_06757_));
 sky130_fd_sc_hd__o21ba_2 _21074_ (.A1(_06626_),
    .A2(_06630_),
    .B1_N(_06628_),
    .X(_06758_));
 sky130_fd_sc_hd__a2bb2o_2 _21075_ (.A1_N(_06757_),
    .A2_N(_06758_),
    .B1(_06757_),
    .B2(_06758_),
    .X(_06759_));
 sky130_fd_sc_hd__a2bb2o_2 _21076_ (.A1_N(_06747_),
    .A2_N(_06759_),
    .B1(_06747_),
    .B2(_06759_),
    .X(_06760_));
 sky130_fd_sc_hd__o22a_2 _21077_ (.A1(_06631_),
    .A2(_06632_),
    .B1(_06622_),
    .B2(_06633_),
    .X(_06761_));
 sky130_fd_sc_hd__a2bb2o_2 _21078_ (.A1_N(_06760_),
    .A2_N(_06761_),
    .B1(_06760_),
    .B2(_06761_),
    .X(_06762_));
 sky130_fd_sc_hd__a2bb2o_2 _21079_ (.A1_N(_06740_),
    .A2_N(_06762_),
    .B1(_06740_),
    .B2(_06762_),
    .X(_06763_));
 sky130_fd_sc_hd__o22a_2 _21080_ (.A1(_06641_),
    .A2(_06646_),
    .B1(_06640_),
    .B2(_06647_),
    .X(_06764_));
 sky130_fd_sc_hd__o22a_2 _21081_ (.A1(_06666_),
    .A2(_06667_),
    .B1(_06661_),
    .B2(_06668_),
    .X(_06765_));
 sky130_fd_sc_hd__o21ba_2 _21082_ (.A1(_06642_),
    .A2(_06645_),
    .B1_N(_06643_),
    .X(_06766_));
 sky130_fd_sc_hd__o21ba_2 _21083_ (.A1(_06657_),
    .A2(_06660_),
    .B1_N(_06658_),
    .X(_06767_));
 sky130_fd_sc_hd__or2_2 _21084_ (.A(_05735_),
    .B(_06502_),
    .X(_06768_));
 sky130_fd_sc_hd__and4_2 _21085_ (.A(_05742_),
    .B(_06239_),
    .C(_05744_),
    .D(_06371_),
    .X(_06769_));
 sky130_fd_sc_hd__o22a_2 _21086_ (.A1(_05738_),
    .A2(_06236_),
    .B1(_05739_),
    .B2(_05986_),
    .X(_06770_));
 sky130_fd_sc_hd__or2_2 _21087_ (.A(_06769_),
    .B(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__a2bb2o_2 _21088_ (.A1_N(_06768_),
    .A2_N(_06771_),
    .B1(_06768_),
    .B2(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__a2bb2o_2 _21089_ (.A1_N(_06767_),
    .A2_N(_06772_),
    .B1(_06767_),
    .B2(_06772_),
    .X(_06773_));
 sky130_fd_sc_hd__a2bb2o_2 _21090_ (.A1_N(_06766_),
    .A2_N(_06773_),
    .B1(_06766_),
    .B2(_06773_),
    .X(_06774_));
 sky130_fd_sc_hd__a2bb2o_2 _21091_ (.A1_N(_06765_),
    .A2_N(_06774_),
    .B1(_06765_),
    .B2(_06774_),
    .X(_06775_));
 sky130_fd_sc_hd__a2bb2o_2 _21092_ (.A1_N(_06764_),
    .A2_N(_06775_),
    .B1(_06764_),
    .B2(_06775_),
    .X(_06776_));
 sky130_fd_sc_hd__o22a_2 _21093_ (.A1(_06639_),
    .A2(_06648_),
    .B1(_06638_),
    .B2(_06649_),
    .X(_06777_));
 sky130_fd_sc_hd__a2bb2o_2 _21094_ (.A1_N(_06776_),
    .A2_N(_06777_),
    .B1(_06776_),
    .B2(_06777_),
    .X(_06778_));
 sky130_fd_sc_hd__a2bb2o_2 _21095_ (.A1_N(_06763_),
    .A2_N(_06778_),
    .B1(_06763_),
    .B2(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__a2bb2o_2 _21096_ (.A1_N(_06739_),
    .A2_N(_06779_),
    .B1(_06739_),
    .B2(_06779_),
    .X(_06780_));
 sky130_fd_sc_hd__a2bb2o_2 _21097_ (.A1_N(_06738_),
    .A2_N(_06780_),
    .B1(_06738_),
    .B2(_06780_),
    .X(_06781_));
 sky130_fd_sc_hd__o22a_2 _21098_ (.A1(_06678_),
    .A2(_06679_),
    .B1(_06669_),
    .B2(_06680_),
    .X(_06782_));
 sky130_fd_sc_hd__o22a_2 _21099_ (.A1(_06566_),
    .A2(_06714_),
    .B1(_06699_),
    .B2(_06715_),
    .X(_06783_));
 sky130_fd_sc_hd__or2_2 _21100_ (.A(_06168_),
    .B(_05815_),
    .X(_06784_));
 sky130_fd_sc_hd__o22a_2 _21101_ (.A1(_06299_),
    .A2(_05509_),
    .B1(_06300_),
    .B2(_05606_),
    .X(_06785_));
 sky130_fd_sc_hd__and4_2 _21102_ (.A(_06171_),
    .B(_11912_),
    .C(_06172_),
    .D(_11910_),
    .X(_06786_));
 sky130_fd_sc_hd__or2_2 _21103_ (.A(_06785_),
    .B(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__a2bb2o_2 _21104_ (.A1_N(_06784_),
    .A2_N(_06787_),
    .B1(_06784_),
    .B2(_06787_),
    .X(_06788_));
 sky130_fd_sc_hd__or2_2 _21105_ (.A(_06176_),
    .B(_05828_),
    .X(_06789_));
 sky130_fd_sc_hd__and4_2 _21106_ (.A(_06182_),
    .B(_11919_),
    .C(_06183_),
    .D(_11916_),
    .X(_06790_));
 sky130_fd_sc_hd__o22a_2 _21107_ (.A1(_06307_),
    .A2(_05255_),
    .B1(_06415_),
    .B2(_06014_),
    .X(_06791_));
 sky130_fd_sc_hd__or2_2 _21108_ (.A(_06790_),
    .B(_06791_),
    .X(_06792_));
 sky130_fd_sc_hd__a2bb2o_2 _21109_ (.A1_N(_06789_),
    .A2_N(_06792_),
    .B1(_06789_),
    .B2(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__o21ba_2 _21110_ (.A1(_06662_),
    .A2(_06665_),
    .B1_N(_06663_),
    .X(_06794_));
 sky130_fd_sc_hd__a2bb2o_2 _21111_ (.A1_N(_06793_),
    .A2_N(_06794_),
    .B1(_06793_),
    .B2(_06794_),
    .X(_06795_));
 sky130_fd_sc_hd__a2bb2o_2 _21112_ (.A1_N(_06788_),
    .A2_N(_06795_),
    .B1(_06788_),
    .B2(_06795_),
    .X(_06796_));
 sky130_fd_sc_hd__o21ba_2 _21113_ (.A1(_06672_),
    .A2(_06675_),
    .B1_N(_06673_),
    .X(_06797_));
 sky130_fd_sc_hd__o21ba_2 _21114_ (.A1(_06701_),
    .A2(_06705_),
    .B1_N(_06704_),
    .X(_06798_));
 sky130_fd_sc_hd__or2_2 _21115_ (.A(_05309_),
    .B(_05736_),
    .X(_06799_));
 sky130_fd_sc_hd__and4_2 _21116_ (.A(_06425_),
    .B(_05743_),
    .C(_06426_),
    .D(_05514_),
    .X(_06800_));
 sky130_fd_sc_hd__o22a_2 _21117_ (.A1(_06428_),
    .A2(_05345_),
    .B1(_05388_),
    .B2(_05157_),
    .X(_06801_));
 sky130_fd_sc_hd__or2_2 _21118_ (.A(_06800_),
    .B(_06801_),
    .X(_06802_));
 sky130_fd_sc_hd__a2bb2o_2 _21119_ (.A1_N(_06799_),
    .A2_N(_06802_),
    .B1(_06799_),
    .B2(_06802_),
    .X(_06803_));
 sky130_fd_sc_hd__a2bb2o_2 _21120_ (.A1_N(_06798_),
    .A2_N(_06803_),
    .B1(_06798_),
    .B2(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__a2bb2o_2 _21121_ (.A1_N(_06797_),
    .A2_N(_06804_),
    .B1(_06797_),
    .B2(_06804_),
    .X(_06805_));
 sky130_fd_sc_hd__o22a_2 _21122_ (.A1(_06671_),
    .A2(_06676_),
    .B1(_06670_),
    .B2(_06677_),
    .X(_06806_));
 sky130_fd_sc_hd__a2bb2o_2 _21123_ (.A1_N(_06805_),
    .A2_N(_06806_),
    .B1(_06805_),
    .B2(_06806_),
    .X(_06807_));
 sky130_fd_sc_hd__a2bb2o_2 _21124_ (.A1_N(_06796_),
    .A2_N(_06807_),
    .B1(_06796_),
    .B2(_06807_),
    .X(_06808_));
 sky130_fd_sc_hd__a2bb2o_2 _21125_ (.A1_N(_06783_),
    .A2_N(_06808_),
    .B1(_06783_),
    .B2(_06808_),
    .X(_06809_));
 sky130_fd_sc_hd__a2bb2o_2 _21126_ (.A1_N(_06782_),
    .A2_N(_06809_),
    .B1(_06782_),
    .B2(_06809_),
    .X(_06810_));
 sky130_fd_sc_hd__o22a_2 _21127_ (.A1(_06711_),
    .A2(_06712_),
    .B1(_06706_),
    .B2(_06713_),
    .X(_06811_));
 sky130_fd_sc_hd__or2_2 _21128_ (.A(_06451_),
    .B(_05164_),
    .X(_06812_));
 sky130_fd_sc_hd__o22a_2 _21129_ (.A1(_06572_),
    .A2(_05172_),
    .B1(_06573_),
    .B2(_06429_),
    .X(_06813_));
 sky130_fd_sc_hd__and4_2 _21130_ (.A(_06453_),
    .B(_05176_),
    .C(_06280_),
    .D(_05781_),
    .X(_06814_));
 sky130_fd_sc_hd__or2_2 _21131_ (.A(_06813_),
    .B(_06814_),
    .X(_06815_));
 sky130_fd_sc_hd__a2bb2o_2 _21132_ (.A1_N(_06812_),
    .A2_N(_06815_),
    .B1(_06812_),
    .B2(_06815_),
    .X(_06816_));
 sky130_fd_sc_hd__or2_2 _21133_ (.A(_05926_),
    .B(_05191_),
    .X(_06817_));
 sky130_fd_sc_hd__buf_1 _21134_ (.A(_06579_),
    .X(_06818_));
 sky130_fd_sc_hd__o22a_2 _21135_ (.A1(_06818_),
    .A2(_05225_),
    .B1(_06030_),
    .B2(_05312_),
    .X(_06819_));
 sky130_fd_sc_hd__and4_2 _21136_ (.A(_11585_),
    .B(_11943_),
    .C(_11589_),
    .D(_05198_),
    .X(_06820_));
 sky130_fd_sc_hd__or2_2 _21137_ (.A(_06819_),
    .B(_06820_),
    .X(_06821_));
 sky130_fd_sc_hd__a2bb2o_2 _21138_ (.A1_N(_06817_),
    .A2_N(_06821_),
    .B1(_06817_),
    .B2(_06821_),
    .X(_06822_));
 sky130_fd_sc_hd__o21ba_2 _21139_ (.A1(_06707_),
    .A2(_06710_),
    .B1_N(_06708_),
    .X(_06823_));
 sky130_fd_sc_hd__a2bb2o_2 _21140_ (.A1_N(_06822_),
    .A2_N(_06823_),
    .B1(_06822_),
    .B2(_06823_),
    .X(_06824_));
 sky130_fd_sc_hd__a2bb2o_2 _21141_ (.A1_N(_06816_),
    .A2_N(_06824_),
    .B1(_06816_),
    .B2(_06824_),
    .X(_06825_));
 sky130_fd_sc_hd__a2bb2o_2 _21142_ (.A1_N(_06695_),
    .A2_N(_06825_),
    .B1(_06695_),
    .B2(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__a2bb2o_2 _21143_ (.A1_N(_06811_),
    .A2_N(_06826_),
    .B1(_06811_),
    .B2(_06826_),
    .X(_06827_));
 sky130_vsdinv _21144_ (.A(\pcpi_mul.rs2[28] ),
    .Y(_06828_));
 sky130_fd_sc_hd__buf_1 _21145_ (.A(_06828_),
    .X(_06829_));
 sky130_fd_sc_hd__buf_1 _21146_ (.A(_06829_),
    .X(_06830_));
 sky130_fd_sc_hd__buf_1 _21147_ (.A(_06830_),
    .X(_06831_));
 sky130_fd_sc_hd__o22a_2 _21148_ (.A1(_06831_),
    .A2(_04544_),
    .B1(_06687_),
    .B2(_04689_),
    .X(_06832_));
 sky130_fd_sc_hd__buf_1 _21149_ (.A(_06829_),
    .X(_06833_));
 sky130_fd_sc_hd__or4_2 _21150_ (.A(_06833_),
    .B(_04543_),
    .C(_06685_),
    .D(_04703_),
    .X(_06834_));
 sky130_fd_sc_hd__or2b_2 _21151_ (.A(_06832_),
    .B_N(_06834_),
    .X(_06835_));
 sky130_fd_sc_hd__o21ba_2 _21152_ (.A1(_06689_),
    .A2(_06692_),
    .B1_N(_06691_),
    .X(_06836_));
 sky130_fd_sc_hd__or2_2 _21153_ (.A(_06271_),
    .B(_05137_),
    .X(_06837_));
 sky130_fd_sc_hd__o22a_2 _21154_ (.A1(_06562_),
    .A2(_04701_),
    .B1(_06440_),
    .B2(_05141_),
    .X(_06838_));
 sky130_fd_sc_hd__and4_2 _21155_ (.A(_11574_),
    .B(_05144_),
    .C(_11579_),
    .D(_11948_),
    .X(_06839_));
 sky130_fd_sc_hd__or2_2 _21156_ (.A(_06838_),
    .B(_06839_),
    .X(_06840_));
 sky130_fd_sc_hd__a2bb2o_2 _21157_ (.A1_N(_06837_),
    .A2_N(_06840_),
    .B1(_06837_),
    .B2(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__or2_2 _21158_ (.A(_06836_),
    .B(_06841_),
    .X(_06842_));
 sky130_fd_sc_hd__a21bo_2 _21159_ (.A1(_06836_),
    .A2(_06841_),
    .B1_N(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__or2_2 _21160_ (.A(_06835_),
    .B(_06843_),
    .X(_06844_));
 sky130_fd_sc_hd__a21bo_2 _21161_ (.A1(_06835_),
    .A2(_06843_),
    .B1_N(_06844_),
    .X(_06845_));
 sky130_fd_sc_hd__a2bb2o_2 _21162_ (.A1_N(_06697_),
    .A2_N(_06845_),
    .B1(_06697_),
    .B2(_06845_),
    .X(_06846_));
 sky130_fd_sc_hd__a2bb2o_2 _21163_ (.A1_N(_06827_),
    .A2_N(_06846_),
    .B1(_06827_),
    .B2(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__a2bb2o_2 _21164_ (.A1_N(_06717_),
    .A2_N(_06847_),
    .B1(_06717_),
    .B2(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__a2bb2o_2 _21165_ (.A1_N(_06810_),
    .A2_N(_06848_),
    .B1(_06810_),
    .B2(_06848_),
    .X(_06849_));
 sky130_fd_sc_hd__o22a_2 _21166_ (.A1(_06589_),
    .A2(_06718_),
    .B1(_06683_),
    .B2(_06719_),
    .X(_06850_));
 sky130_fd_sc_hd__a2bb2o_2 _21167_ (.A1_N(_06849_),
    .A2_N(_06850_),
    .B1(_06849_),
    .B2(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__a2bb2o_2 _21168_ (.A1_N(_06781_),
    .A2_N(_06851_),
    .B1(_06781_),
    .B2(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__o22a_2 _21169_ (.A1(_06720_),
    .A2(_06721_),
    .B1(_06655_),
    .B2(_06722_),
    .X(_06853_));
 sky130_fd_sc_hd__a2bb2o_2 _21170_ (.A1_N(_06852_),
    .A2_N(_06853_),
    .B1(_06852_),
    .B2(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__a2bb2o_2 _21171_ (.A1_N(_06737_),
    .A2_N(_06854_),
    .B1(_06737_),
    .B2(_06854_),
    .X(_06855_));
 sky130_fd_sc_hd__o22a_2 _21172_ (.A1(_06723_),
    .A2(_06724_),
    .B1(_06611_),
    .B2(_06725_),
    .X(_06856_));
 sky130_fd_sc_hd__a2bb2o_2 _21173_ (.A1_N(_06855_),
    .A2_N(_06856_),
    .B1(_06855_),
    .B2(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__a2bb2o_2 _21174_ (.A1_N(_06610_),
    .A2_N(_06857_),
    .B1(_06610_),
    .B2(_06857_),
    .X(_06858_));
 sky130_fd_sc_hd__o22a_2 _21175_ (.A1(_06726_),
    .A2(_06727_),
    .B1(_06485_),
    .B2(_06728_),
    .X(_06859_));
 sky130_fd_sc_hd__or2_2 _21176_ (.A(_06858_),
    .B(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__a21bo_2 _21177_ (.A1(_06858_),
    .A2(_06859_),
    .B1_N(_06860_),
    .X(_06861_));
 sky130_fd_sc_hd__or2_2 _21178_ (.A(_06604_),
    .B(_06732_),
    .X(_06862_));
 sky130_fd_sc_hd__or3_2 _21179_ (.A(_06342_),
    .B(_06481_),
    .C(_06862_),
    .X(_06863_));
 sky130_fd_sc_hd__o221a_2 _21180_ (.A1(_06603_),
    .A2(_06730_),
    .B1(_06605_),
    .B2(_06862_),
    .C1(_06731_),
    .X(_06864_));
 sky130_fd_sc_hd__o21ai_2 _21181_ (.A1(_06349_),
    .A2(_06863_),
    .B1(_06864_),
    .Y(_06865_));
 sky130_vsdinv _21182_ (.A(_06865_),
    .Y(_06866_));
 sky130_vsdinv _21183_ (.A(_06861_),
    .Y(_06867_));
 sky130_fd_sc_hd__o22a_2 _21184_ (.A1(_06861_),
    .A2(_06866_),
    .B1(_06867_),
    .B2(_06865_),
    .X(_02647_));
 sky130_fd_sc_hd__o22a_2 _21185_ (.A1(_06855_),
    .A2(_06856_),
    .B1(_06610_),
    .B2(_06857_),
    .X(_06868_));
 sky130_fd_sc_hd__o22a_2 _21186_ (.A1(_06739_),
    .A2(_06779_),
    .B1(_06738_),
    .B2(_06780_),
    .X(_06869_));
 sky130_fd_sc_hd__o22a_2 _21187_ (.A1(_06760_),
    .A2(_06761_),
    .B1(_06740_),
    .B2(_06762_),
    .X(_06870_));
 sky130_fd_sc_hd__or2_2 _21188_ (.A(_06869_),
    .B(_06870_),
    .X(_06871_));
 sky130_fd_sc_hd__a21bo_2 _21189_ (.A1(_06869_),
    .A2(_06870_),
    .B1_N(_06871_),
    .X(_06872_));
 sky130_fd_sc_hd__o22a_2 _21190_ (.A1(_06776_),
    .A2(_06777_),
    .B1(_06763_),
    .B2(_06778_),
    .X(_06873_));
 sky130_fd_sc_hd__o22a_2 _21191_ (.A1(_06783_),
    .A2(_06808_),
    .B1(_06782_),
    .B2(_06809_),
    .X(_06874_));
 sky130_fd_sc_hd__o21ba_2 _21192_ (.A1(_06745_),
    .A2(_06746_),
    .B1_N(_06741_),
    .X(_06875_));
 sky130_fd_sc_hd__buf_1 _21193_ (.A(_11882_),
    .X(_06876_));
 sky130_fd_sc_hd__and4_2 _21194_ (.A(_11637_),
    .B(_11885_),
    .C(_11643_),
    .D(_06876_),
    .X(_06877_));
 sky130_fd_sc_hd__buf_1 _21195_ (.A(_06623_),
    .X(_06878_));
 sky130_fd_sc_hd__buf_1 _21196_ (.A(_06878_),
    .X(_06879_));
 sky130_fd_sc_hd__o22a_2 _21197_ (.A1(_05153_),
    .A2(_06879_),
    .B1(_05156_),
    .B2(_06750_),
    .X(_06880_));
 sky130_fd_sc_hd__or2_2 _21198_ (.A(_06877_),
    .B(_06880_),
    .X(_06881_));
 sky130_fd_sc_hd__buf_1 _21199_ (.A(_06496_),
    .X(_06882_));
 sky130_fd_sc_hd__or2_2 _21200_ (.A(_05162_),
    .B(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__a2bb2o_2 _21201_ (.A1_N(_06881_),
    .A2_N(_06883_),
    .B1(_06881_),
    .B2(_06883_),
    .X(_06884_));
 sky130_fd_sc_hd__buf_1 _21202_ (.A(\pcpi_mul.rs1[25] ),
    .X(_06885_));
 sky130_fd_sc_hd__and4_2 _21203_ (.A(_11628_),
    .B(_06752_),
    .C(_11632_),
    .D(_06885_),
    .X(_06886_));
 sky130_fd_sc_hd__o22a_2 _21204_ (.A1(_05826_),
    .A2(_06233_),
    .B1(_05827_),
    .B2(_06616_),
    .X(_06887_));
 sky130_fd_sc_hd__or2_2 _21205_ (.A(_06886_),
    .B(_06887_),
    .X(_06888_));
 sky130_vsdinv _21206_ (.A(\pcpi_mul.rs1[29] ),
    .Y(_06889_));
 sky130_fd_sc_hd__buf_1 _21207_ (.A(_06889_),
    .X(_06890_));
 sky130_fd_sc_hd__buf_1 _21208_ (.A(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__or2_2 _21209_ (.A(_05713_),
    .B(_06891_),
    .X(_06892_));
 sky130_fd_sc_hd__a2bb2o_2 _21210_ (.A1_N(_06888_),
    .A2_N(_06892_),
    .B1(_06888_),
    .B2(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__o21ba_2 _21211_ (.A1(_06751_),
    .A2(_06756_),
    .B1_N(_06753_),
    .X(_06894_));
 sky130_fd_sc_hd__a2bb2o_2 _21212_ (.A1_N(_06893_),
    .A2_N(_06894_),
    .B1(_06893_),
    .B2(_06894_),
    .X(_06895_));
 sky130_fd_sc_hd__a2bb2o_2 _21213_ (.A1_N(_06884_),
    .A2_N(_06895_),
    .B1(_06884_),
    .B2(_06895_),
    .X(_06896_));
 sky130_fd_sc_hd__o22a_2 _21214_ (.A1(_06757_),
    .A2(_06758_),
    .B1(_06747_),
    .B2(_06759_),
    .X(_06897_));
 sky130_fd_sc_hd__a2bb2o_2 _21215_ (.A1_N(_06896_),
    .A2_N(_06897_),
    .B1(_06896_),
    .B2(_06897_),
    .X(_06898_));
 sky130_fd_sc_hd__a2bb2o_2 _21216_ (.A1_N(_06875_),
    .A2_N(_06898_),
    .B1(_06875_),
    .B2(_06898_),
    .X(_06899_));
 sky130_fd_sc_hd__o22a_2 _21217_ (.A1(_06767_),
    .A2(_06772_),
    .B1(_06766_),
    .B2(_06773_),
    .X(_06900_));
 sky130_fd_sc_hd__o22a_2 _21218_ (.A1(_06793_),
    .A2(_06794_),
    .B1(_06788_),
    .B2(_06795_),
    .X(_06901_));
 sky130_fd_sc_hd__o21ba_2 _21219_ (.A1(_06768_),
    .A2(_06771_),
    .B1_N(_06769_),
    .X(_06902_));
 sky130_fd_sc_hd__o21ba_2 _21220_ (.A1(_06784_),
    .A2(_06787_),
    .B1_N(_06786_),
    .X(_06903_));
 sky130_fd_sc_hd__buf_1 _21221_ (.A(_05994_),
    .X(_06904_));
 sky130_fd_sc_hd__o22a_2 _21222_ (.A1(_06132_),
    .A2(_06501_),
    .B1(_04828_),
    .B2(_06904_),
    .X(_06905_));
 sky130_fd_sc_hd__and4_2 _21223_ (.A(_11620_),
    .B(_06371_),
    .C(_11624_),
    .D(_11899_),
    .X(_06906_));
 sky130_fd_sc_hd__nor2_2 _21224_ (.A(_06905_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__nor2_2 _21225_ (.A(_04795_),
    .B(_06112_),
    .Y(_06908_));
 sky130_fd_sc_hd__a2bb2o_2 _21226_ (.A1_N(_06907_),
    .A2_N(_06908_),
    .B1(_06907_),
    .B2(_06908_),
    .X(_06909_));
 sky130_fd_sc_hd__a2bb2o_2 _21227_ (.A1_N(_06903_),
    .A2_N(_06909_),
    .B1(_06903_),
    .B2(_06909_),
    .X(_06910_));
 sky130_fd_sc_hd__a2bb2o_2 _21228_ (.A1_N(_06902_),
    .A2_N(_06910_),
    .B1(_06902_),
    .B2(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__a2bb2o_2 _21229_ (.A1_N(_06901_),
    .A2_N(_06911_),
    .B1(_06901_),
    .B2(_06911_),
    .X(_06912_));
 sky130_fd_sc_hd__a2bb2o_2 _21230_ (.A1_N(_06900_),
    .A2_N(_06912_),
    .B1(_06900_),
    .B2(_06912_),
    .X(_06913_));
 sky130_fd_sc_hd__o22a_2 _21231_ (.A1(_06765_),
    .A2(_06774_),
    .B1(_06764_),
    .B2(_06775_),
    .X(_06914_));
 sky130_fd_sc_hd__a2bb2o_2 _21232_ (.A1_N(_06913_),
    .A2_N(_06914_),
    .B1(_06913_),
    .B2(_06914_),
    .X(_06915_));
 sky130_fd_sc_hd__a2bb2o_2 _21233_ (.A1_N(_06899_),
    .A2_N(_06915_),
    .B1(_06899_),
    .B2(_06915_),
    .X(_06916_));
 sky130_fd_sc_hd__a2bb2o_2 _21234_ (.A1_N(_06874_),
    .A2_N(_06916_),
    .B1(_06874_),
    .B2(_06916_),
    .X(_06917_));
 sky130_fd_sc_hd__a2bb2o_2 _21235_ (.A1_N(_06873_),
    .A2_N(_06917_),
    .B1(_06873_),
    .B2(_06917_),
    .X(_06918_));
 sky130_fd_sc_hd__o22a_2 _21236_ (.A1(_06805_),
    .A2(_06806_),
    .B1(_06796_),
    .B2(_06807_),
    .X(_06919_));
 sky130_fd_sc_hd__o22a_2 _21237_ (.A1(_06695_),
    .A2(_06825_),
    .B1(_06811_),
    .B2(_06826_),
    .X(_06920_));
 sky130_fd_sc_hd__or2_2 _21238_ (.A(_06168_),
    .B(_06237_),
    .X(_06921_));
 sky130_fd_sc_hd__o22a_2 _21239_ (.A1(_06299_),
    .A2(_05606_),
    .B1(_06300_),
    .B2(_05814_),
    .X(_06922_));
 sky130_fd_sc_hd__and4_2 _21240_ (.A(_06171_),
    .B(_11910_),
    .C(_06172_),
    .D(_06517_),
    .X(_06923_));
 sky130_fd_sc_hd__or2_2 _21241_ (.A(_06922_),
    .B(_06923_),
    .X(_06924_));
 sky130_fd_sc_hd__a2bb2o_2 _21242_ (.A1_N(_06921_),
    .A2_N(_06924_),
    .B1(_06921_),
    .B2(_06924_),
    .X(_06925_));
 sky130_fd_sc_hd__or2_2 _21243_ (.A(_06176_),
    .B(_05895_),
    .X(_06926_));
 sky130_fd_sc_hd__o22a_2 _21244_ (.A1(_05945_),
    .A2(_05342_),
    .B1(_06415_),
    .B2(_05428_),
    .X(_06927_));
 sky130_fd_sc_hd__buf_1 _21245_ (.A(\pcpi_mul.rs2[14] ),
    .X(_06928_));
 sky130_fd_sc_hd__buf_1 _21246_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06929_));
 sky130_fd_sc_hd__and4_2 _21247_ (.A(_06928_),
    .B(_11916_),
    .C(_06929_),
    .D(_11914_),
    .X(_06930_));
 sky130_fd_sc_hd__or2_2 _21248_ (.A(_06927_),
    .B(_06930_),
    .X(_06931_));
 sky130_fd_sc_hd__a2bb2o_2 _21249_ (.A1_N(_06926_),
    .A2_N(_06931_),
    .B1(_06926_),
    .B2(_06931_),
    .X(_06932_));
 sky130_fd_sc_hd__o21ba_2 _21250_ (.A1(_06789_),
    .A2(_06792_),
    .B1_N(_06790_),
    .X(_06933_));
 sky130_fd_sc_hd__a2bb2o_2 _21251_ (.A1_N(_06932_),
    .A2_N(_06933_),
    .B1(_06932_),
    .B2(_06933_),
    .X(_06934_));
 sky130_fd_sc_hd__a2bb2o_2 _21252_ (.A1_N(_06925_),
    .A2_N(_06934_),
    .B1(_06925_),
    .B2(_06934_),
    .X(_06935_));
 sky130_fd_sc_hd__o21ba_2 _21253_ (.A1(_06799_),
    .A2(_06802_),
    .B1_N(_06800_),
    .X(_06936_));
 sky130_fd_sc_hd__o21ba_2 _21254_ (.A1(_06812_),
    .A2(_06815_),
    .B1_N(_06814_),
    .X(_06937_));
 sky130_fd_sc_hd__or2_2 _21255_ (.A(_05393_),
    .B(_05845_),
    .X(_06938_));
 sky130_fd_sc_hd__o22a_2 _21256_ (.A1(_06428_),
    .A2(_05431_),
    .B1(_06549_),
    .B2(_05609_),
    .X(_06939_));
 sky130_fd_sc_hd__and4_2 _21257_ (.A(_06425_),
    .B(_05514_),
    .C(_06426_),
    .D(_05516_),
    .X(_06940_));
 sky130_fd_sc_hd__or2_2 _21258_ (.A(_06939_),
    .B(_06940_),
    .X(_06941_));
 sky130_fd_sc_hd__a2bb2o_2 _21259_ (.A1_N(_06938_),
    .A2_N(_06941_),
    .B1(_06938_),
    .B2(_06941_),
    .X(_06942_));
 sky130_fd_sc_hd__a2bb2o_2 _21260_ (.A1_N(_06937_),
    .A2_N(_06942_),
    .B1(_06937_),
    .B2(_06942_),
    .X(_06943_));
 sky130_fd_sc_hd__a2bb2o_2 _21261_ (.A1_N(_06936_),
    .A2_N(_06943_),
    .B1(_06936_),
    .B2(_06943_),
    .X(_06944_));
 sky130_fd_sc_hd__o22a_2 _21262_ (.A1(_06798_),
    .A2(_06803_),
    .B1(_06797_),
    .B2(_06804_),
    .X(_06945_));
 sky130_fd_sc_hd__a2bb2o_2 _21263_ (.A1_N(_06944_),
    .A2_N(_06945_),
    .B1(_06944_),
    .B2(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__a2bb2o_2 _21264_ (.A1_N(_06935_),
    .A2_N(_06946_),
    .B1(_06935_),
    .B2(_06946_),
    .X(_06947_));
 sky130_fd_sc_hd__a2bb2o_2 _21265_ (.A1_N(_06920_),
    .A2_N(_06947_),
    .B1(_06920_),
    .B2(_06947_),
    .X(_06948_));
 sky130_fd_sc_hd__a2bb2o_2 _21266_ (.A1_N(_06919_),
    .A2_N(_06948_),
    .B1(_06919_),
    .B2(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__o22a_2 _21267_ (.A1(_06822_),
    .A2(_06823_),
    .B1(_06816_),
    .B2(_06824_),
    .X(_06950_));
 sky130_fd_sc_hd__or2_2 _21268_ (.A(_06451_),
    .B(_05072_),
    .X(_06951_));
 sky130_fd_sc_hd__o22a_2 _21269_ (.A1(_06572_),
    .A2(_05076_),
    .B1(_06573_),
    .B2(_05258_),
    .X(_06952_));
 sky130_fd_sc_hd__and4_2 _21270_ (.A(_06453_),
    .B(_05177_),
    .C(_06280_),
    .D(_05260_),
    .X(_06953_));
 sky130_fd_sc_hd__or2_2 _21271_ (.A(_06952_),
    .B(_06953_),
    .X(_06954_));
 sky130_fd_sc_hd__a2bb2o_2 _21272_ (.A1_N(_06951_),
    .A2_N(_06954_),
    .B1(_06951_),
    .B2(_06954_),
    .X(_06955_));
 sky130_fd_sc_hd__or2_2 _21273_ (.A(_06035_),
    .B(_06568_),
    .X(_06956_));
 sky130_fd_sc_hd__o22a_2 _21274_ (.A1(_06818_),
    .A2(_05195_),
    .B1(_06033_),
    .B2(_05575_),
    .X(_06957_));
 sky130_fd_sc_hd__and4_2 _21275_ (.A(_11585_),
    .B(_05198_),
    .C(_11589_),
    .D(_05577_),
    .X(_06958_));
 sky130_fd_sc_hd__or2_2 _21276_ (.A(_06957_),
    .B(_06958_),
    .X(_06959_));
 sky130_fd_sc_hd__a2bb2o_2 _21277_ (.A1_N(_06956_),
    .A2_N(_06959_),
    .B1(_06956_),
    .B2(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__o21ba_2 _21278_ (.A1(_06817_),
    .A2(_06821_),
    .B1_N(_06820_),
    .X(_06961_));
 sky130_fd_sc_hd__a2bb2o_2 _21279_ (.A1_N(_06960_),
    .A2_N(_06961_),
    .B1(_06960_),
    .B2(_06961_),
    .X(_06962_));
 sky130_fd_sc_hd__a2bb2o_2 _21280_ (.A1_N(_06955_),
    .A2_N(_06962_),
    .B1(_06955_),
    .B2(_06962_),
    .X(_06963_));
 sky130_fd_sc_hd__a2bb2o_2 _21281_ (.A1_N(_06842_),
    .A2_N(_06963_),
    .B1(_06842_),
    .B2(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__a2bb2o_2 _21282_ (.A1_N(_06950_),
    .A2_N(_06964_),
    .B1(_06950_),
    .B2(_06964_),
    .X(_06965_));
 sky130_fd_sc_hd__or2_2 _21283_ (.A(_06684_),
    .B(_04702_),
    .X(_06966_));
 sky130_fd_sc_hd__and4_2 _21284_ (.A(_11570_),
    .B(_11955_),
    .C(\pcpi_mul.rs2[29] ),
    .D(_11957_),
    .X(_06967_));
 sky130_vsdinv _21285_ (.A(\pcpi_mul.rs2[29] ),
    .Y(_06968_));
 sky130_fd_sc_hd__o22a_2 _21286_ (.A1(_06828_),
    .A2(_04709_),
    .B1(_06968_),
    .B2(_04710_),
    .X(_06969_));
 sky130_fd_sc_hd__or2_2 _21287_ (.A(_06967_),
    .B(_06969_),
    .X(_06970_));
 sky130_fd_sc_hd__a2bb2o_2 _21288_ (.A1_N(_06966_),
    .A2_N(_06970_),
    .B1(_06966_),
    .B2(_06970_),
    .X(_06971_));
 sky130_fd_sc_hd__o21ba_2 _21289_ (.A1(_06837_),
    .A2(_06840_),
    .B1_N(_06839_),
    .X(_06972_));
 sky130_fd_sc_hd__or2_2 _21290_ (.A(_06272_),
    .B(_06151_),
    .X(_06973_));
 sky130_fd_sc_hd__buf_1 _21291_ (.A(_06562_),
    .X(_06974_));
 sky130_fd_sc_hd__o22a_2 _21292_ (.A1(_06974_),
    .A2(_05141_),
    .B1(_06441_),
    .B2(_05227_),
    .X(_06975_));
 sky130_fd_sc_hd__and4_2 _21293_ (.A(_11574_),
    .B(_11949_),
    .C(_11579_),
    .D(_05316_),
    .X(_06976_));
 sky130_fd_sc_hd__or2_2 _21294_ (.A(_06975_),
    .B(_06976_),
    .X(_06977_));
 sky130_fd_sc_hd__a2bb2o_2 _21295_ (.A1_N(_06973_),
    .A2_N(_06977_),
    .B1(_06973_),
    .B2(_06977_),
    .X(_06978_));
 sky130_fd_sc_hd__a2bb2o_2 _21296_ (.A1_N(_06834_),
    .A2_N(_06978_),
    .B1(_06834_),
    .B2(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__a2bb2o_2 _21297_ (.A1_N(_06972_),
    .A2_N(_06979_),
    .B1(_06972_),
    .B2(_06979_),
    .X(_06980_));
 sky130_fd_sc_hd__or2_2 _21298_ (.A(_06971_),
    .B(_06980_),
    .X(_06981_));
 sky130_fd_sc_hd__a21bo_2 _21299_ (.A1(_06971_),
    .A2(_06980_),
    .B1_N(_06981_),
    .X(_06982_));
 sky130_fd_sc_hd__a2bb2o_2 _21300_ (.A1_N(_06844_),
    .A2_N(_06982_),
    .B1(_06844_),
    .B2(_06982_),
    .X(_06983_));
 sky130_fd_sc_hd__a2bb2o_2 _21301_ (.A1_N(_06965_),
    .A2_N(_06983_),
    .B1(_06965_),
    .B2(_06983_),
    .X(_06984_));
 sky130_fd_sc_hd__o22a_2 _21302_ (.A1(_06697_),
    .A2(_06845_),
    .B1(_06827_),
    .B2(_06846_),
    .X(_06985_));
 sky130_fd_sc_hd__a2bb2o_2 _21303_ (.A1_N(_06984_),
    .A2_N(_06985_),
    .B1(_06984_),
    .B2(_06985_),
    .X(_06986_));
 sky130_fd_sc_hd__a2bb2o_2 _21304_ (.A1_N(_06949_),
    .A2_N(_06986_),
    .B1(_06949_),
    .B2(_06986_),
    .X(_06987_));
 sky130_fd_sc_hd__o22a_2 _21305_ (.A1(_06717_),
    .A2(_06847_),
    .B1(_06810_),
    .B2(_06848_),
    .X(_06988_));
 sky130_fd_sc_hd__a2bb2o_2 _21306_ (.A1_N(_06987_),
    .A2_N(_06988_),
    .B1(_06987_),
    .B2(_06988_),
    .X(_06989_));
 sky130_fd_sc_hd__a2bb2o_2 _21307_ (.A1_N(_06918_),
    .A2_N(_06989_),
    .B1(_06918_),
    .B2(_06989_),
    .X(_06990_));
 sky130_fd_sc_hd__o22a_2 _21308_ (.A1(_06849_),
    .A2(_06850_),
    .B1(_06781_),
    .B2(_06851_),
    .X(_06991_));
 sky130_fd_sc_hd__a2bb2o_2 _21309_ (.A1_N(_06990_),
    .A2_N(_06991_),
    .B1(_06990_),
    .B2(_06991_),
    .X(_06992_));
 sky130_fd_sc_hd__a2bb2o_2 _21310_ (.A1_N(_06872_),
    .A2_N(_06992_),
    .B1(_06872_),
    .B2(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__o22a_2 _21311_ (.A1(_06852_),
    .A2(_06853_),
    .B1(_06737_),
    .B2(_06854_),
    .X(_06994_));
 sky130_fd_sc_hd__a2bb2o_2 _21312_ (.A1_N(_06993_),
    .A2_N(_06994_),
    .B1(_06993_),
    .B2(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__a2bb2o_2 _21313_ (.A1_N(_06736_),
    .A2_N(_06995_),
    .B1(_06736_),
    .B2(_06995_),
    .X(_06996_));
 sky130_fd_sc_hd__or2_2 _21314_ (.A(_06868_),
    .B(_06996_),
    .X(_06997_));
 sky130_fd_sc_hd__a21bo_2 _21315_ (.A1(_06868_),
    .A2(_06996_),
    .B1_N(_06997_),
    .X(_06998_));
 sky130_fd_sc_hd__o21ai_2 _21316_ (.A1(_06861_),
    .A2(_06866_),
    .B1(_06860_),
    .Y(_06999_));
 sky130_fd_sc_hd__a2bb2o_2 _21317_ (.A1_N(_06998_),
    .A2_N(_06999_),
    .B1(_06998_),
    .B2(_06999_),
    .X(_02648_));
 sky130_fd_sc_hd__o22a_2 _21318_ (.A1(_06874_),
    .A2(_06916_),
    .B1(_06873_),
    .B2(_06917_),
    .X(_07000_));
 sky130_fd_sc_hd__o22a_2 _21319_ (.A1(_06896_),
    .A2(_06897_),
    .B1(_06875_),
    .B2(_06898_),
    .X(_07001_));
 sky130_fd_sc_hd__or2_2 _21320_ (.A(_07000_),
    .B(_07001_),
    .X(_07002_));
 sky130_fd_sc_hd__a21bo_2 _21321_ (.A1(_07000_),
    .A2(_07001_),
    .B1_N(_07002_),
    .X(_07003_));
 sky130_fd_sc_hd__o22a_2 _21322_ (.A1(_06913_),
    .A2(_06914_),
    .B1(_06899_),
    .B2(_06915_),
    .X(_07004_));
 sky130_fd_sc_hd__o22a_2 _21323_ (.A1(_06920_),
    .A2(_06947_),
    .B1(_06919_),
    .B2(_06948_),
    .X(_07005_));
 sky130_fd_sc_hd__o21ba_2 _21324_ (.A1(_06881_),
    .A2(_06883_),
    .B1_N(_06877_),
    .X(_07006_));
 sky130_fd_sc_hd__buf_1 _21325_ (.A(_06749_),
    .X(_07007_));
 sky130_fd_sc_hd__buf_1 _21326_ (.A(_07007_),
    .X(_07008_));
 sky130_fd_sc_hd__buf_1 _21327_ (.A(_06889_),
    .X(_07009_));
 sky130_fd_sc_hd__buf_1 _21328_ (.A(_07009_),
    .X(_07010_));
 sky130_fd_sc_hd__o22a_2 _21329_ (.A1(_05702_),
    .A2(_07008_),
    .B1(_05703_),
    .B2(_07010_),
    .X(_07011_));
 sky130_fd_sc_hd__buf_1 _21330_ (.A(_11880_),
    .X(_07012_));
 sky130_fd_sc_hd__and4_2 _21331_ (.A(_11638_),
    .B(_06876_),
    .C(_11644_),
    .D(_07012_),
    .X(_07013_));
 sky130_fd_sc_hd__nor2_2 _21332_ (.A(_07011_),
    .B(_07013_),
    .Y(_07014_));
 sky130_fd_sc_hd__buf_1 _21333_ (.A(_06879_),
    .X(_07015_));
 sky130_fd_sc_hd__nor2_2 _21334_ (.A(_06107_),
    .B(_07015_),
    .Y(_07016_));
 sky130_fd_sc_hd__a2bb2o_2 _21335_ (.A1_N(_07014_),
    .A2_N(_07016_),
    .B1(_07014_),
    .B2(_07016_),
    .X(_07017_));
 sky130_fd_sc_hd__o22a_2 _21336_ (.A1(_06368_),
    .A2(_06377_),
    .B1(_06369_),
    .B2(_06743_),
    .X(_07018_));
 sky130_fd_sc_hd__and4_2 _21337_ (.A(_11629_),
    .B(_11893_),
    .C(_11633_),
    .D(_11888_),
    .X(_07019_));
 sky130_fd_sc_hd__nor2_2 _21338_ (.A(_07018_),
    .B(_07019_),
    .Y(_07020_));
 sky130_vsdinv _21339_ (.A(\pcpi_mul.rs1[30] ),
    .Y(_07021_));
 sky130_fd_sc_hd__buf_1 _21340_ (.A(_07021_),
    .X(_07022_));
 sky130_fd_sc_hd__buf_1 _21341_ (.A(_07022_),
    .X(_07023_));
 sky130_fd_sc_hd__buf_1 _21342_ (.A(_07023_),
    .X(_07024_));
 sky130_fd_sc_hd__nor2_2 _21343_ (.A(_04538_),
    .B(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__a2bb2o_2 _21344_ (.A1_N(_07020_),
    .A2_N(_07025_),
    .B1(_07020_),
    .B2(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__o21ba_2 _21345_ (.A1(_06888_),
    .A2(_06892_),
    .B1_N(_06886_),
    .X(_07027_));
 sky130_fd_sc_hd__a2bb2o_2 _21346_ (.A1_N(_07026_),
    .A2_N(_07027_),
    .B1(_07026_),
    .B2(_07027_),
    .X(_07028_));
 sky130_fd_sc_hd__a2bb2o_2 _21347_ (.A1_N(_07017_),
    .A2_N(_07028_),
    .B1(_07017_),
    .B2(_07028_),
    .X(_07029_));
 sky130_fd_sc_hd__o22a_2 _21348_ (.A1(_06893_),
    .A2(_06894_),
    .B1(_06884_),
    .B2(_06895_),
    .X(_07030_));
 sky130_fd_sc_hd__a2bb2o_2 _21349_ (.A1_N(_07029_),
    .A2_N(_07030_),
    .B1(_07029_),
    .B2(_07030_),
    .X(_07031_));
 sky130_fd_sc_hd__a2bb2o_2 _21350_ (.A1_N(_07006_),
    .A2_N(_07031_),
    .B1(_07006_),
    .B2(_07031_),
    .X(_07032_));
 sky130_fd_sc_hd__o22a_2 _21351_ (.A1(_06903_),
    .A2(_06909_),
    .B1(_06902_),
    .B2(_06910_),
    .X(_07033_));
 sky130_fd_sc_hd__o22a_2 _21352_ (.A1(_06932_),
    .A2(_06933_),
    .B1(_06925_),
    .B2(_06934_),
    .X(_07034_));
 sky130_fd_sc_hd__a21oi_2 _21353_ (.A1(_06907_),
    .A2(_06908_),
    .B1(_06906_),
    .Y(_07035_));
 sky130_fd_sc_hd__o21ba_2 _21354_ (.A1(_06921_),
    .A2(_06924_),
    .B1_N(_06923_),
    .X(_07036_));
 sky130_fd_sc_hd__o22a_2 _21355_ (.A1(_06132_),
    .A2(_05995_),
    .B1(_06133_),
    .B2(_06754_),
    .X(_07037_));
 sky130_fd_sc_hd__buf_1 _21356_ (.A(\pcpi_mul.rs1[23] ),
    .X(_07038_));
 sky130_fd_sc_hd__and4_2 _21357_ (.A(_06136_),
    .B(_11899_),
    .C(_06137_),
    .D(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__nor2_2 _21358_ (.A(_07037_),
    .B(_07039_),
    .Y(_07040_));
 sky130_fd_sc_hd__nor2_2 _21359_ (.A(_04830_),
    .B(_06234_),
    .Y(_07041_));
 sky130_fd_sc_hd__a2bb2o_2 _21360_ (.A1_N(_07040_),
    .A2_N(_07041_),
    .B1(_07040_),
    .B2(_07041_),
    .X(_07042_));
 sky130_fd_sc_hd__a2bb2o_2 _21361_ (.A1_N(_07036_),
    .A2_N(_07042_),
    .B1(_07036_),
    .B2(_07042_),
    .X(_07043_));
 sky130_fd_sc_hd__a2bb2o_2 _21362_ (.A1_N(_07035_),
    .A2_N(_07043_),
    .B1(_07035_),
    .B2(_07043_),
    .X(_07044_));
 sky130_fd_sc_hd__a2bb2o_2 _21363_ (.A1_N(_07034_),
    .A2_N(_07044_),
    .B1(_07034_),
    .B2(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__a2bb2o_2 _21364_ (.A1_N(_07033_),
    .A2_N(_07045_),
    .B1(_07033_),
    .B2(_07045_),
    .X(_07046_));
 sky130_fd_sc_hd__o22a_2 _21365_ (.A1(_06901_),
    .A2(_06911_),
    .B1(_06900_),
    .B2(_06912_),
    .X(_07047_));
 sky130_fd_sc_hd__a2bb2o_2 _21366_ (.A1_N(_07046_),
    .A2_N(_07047_),
    .B1(_07046_),
    .B2(_07047_),
    .X(_07048_));
 sky130_fd_sc_hd__a2bb2o_2 _21367_ (.A1_N(_07032_),
    .A2_N(_07048_),
    .B1(_07032_),
    .B2(_07048_),
    .X(_07049_));
 sky130_fd_sc_hd__a2bb2o_2 _21368_ (.A1_N(_07005_),
    .A2_N(_07049_),
    .B1(_07005_),
    .B2(_07049_),
    .X(_07050_));
 sky130_fd_sc_hd__a2bb2o_2 _21369_ (.A1_N(_07004_),
    .A2_N(_07050_),
    .B1(_07004_),
    .B2(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__o22a_2 _21370_ (.A1(_06944_),
    .A2(_06945_),
    .B1(_06935_),
    .B2(_06946_),
    .X(_07052_));
 sky130_fd_sc_hd__o22a_2 _21371_ (.A1(_06842_),
    .A2(_06963_),
    .B1(_06950_),
    .B2(_06964_),
    .X(_07053_));
 sky130_fd_sc_hd__or2_2 _21372_ (.A(_05665_),
    .B(_05892_),
    .X(_07054_));
 sky130_fd_sc_hd__o22a_2 _21373_ (.A1(_05779_),
    .A2(_05814_),
    .B1(_05667_),
    .B2(_06236_),
    .X(_07055_));
 sky130_fd_sc_hd__and4_2 _21374_ (.A(_05669_),
    .B(_06517_),
    .C(_05670_),
    .D(_06239_),
    .X(_07056_));
 sky130_fd_sc_hd__or2_2 _21375_ (.A(_07055_),
    .B(_07056_),
    .X(_07057_));
 sky130_fd_sc_hd__a2bb2o_2 _21376_ (.A1_N(_07054_),
    .A2_N(_07057_),
    .B1(_07054_),
    .B2(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__buf_1 _21377_ (.A(_05605_),
    .X(_07059_));
 sky130_fd_sc_hd__or2_2 _21378_ (.A(_06176_),
    .B(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__o22a_2 _21379_ (.A1(_05945_),
    .A2(_05428_),
    .B1(_06415_),
    .B2(_05509_),
    .X(_07061_));
 sky130_fd_sc_hd__and4_2 _21380_ (.A(_06928_),
    .B(_11914_),
    .C(_06929_),
    .D(_11912_),
    .X(_07062_));
 sky130_fd_sc_hd__or2_2 _21381_ (.A(_07061_),
    .B(_07062_),
    .X(_07063_));
 sky130_fd_sc_hd__a2bb2o_2 _21382_ (.A1_N(_07060_),
    .A2_N(_07063_),
    .B1(_07060_),
    .B2(_07063_),
    .X(_07064_));
 sky130_fd_sc_hd__o21ba_2 _21383_ (.A1(_06926_),
    .A2(_06931_),
    .B1_N(_06930_),
    .X(_07065_));
 sky130_fd_sc_hd__a2bb2o_2 _21384_ (.A1_N(_07064_),
    .A2_N(_07065_),
    .B1(_07064_),
    .B2(_07065_),
    .X(_07066_));
 sky130_fd_sc_hd__a2bb2o_2 _21385_ (.A1_N(_07058_),
    .A2_N(_07066_),
    .B1(_07058_),
    .B2(_07066_),
    .X(_07067_));
 sky130_fd_sc_hd__o21ba_2 _21386_ (.A1(_06938_),
    .A2(_06941_),
    .B1_N(_06940_),
    .X(_07068_));
 sky130_fd_sc_hd__o21ba_2 _21387_ (.A1(_06951_),
    .A2(_06954_),
    .B1_N(_06953_),
    .X(_07069_));
 sky130_fd_sc_hd__or2_2 _21388_ (.A(_05393_),
    .B(_05343_),
    .X(_07070_));
 sky130_fd_sc_hd__o22a_2 _21389_ (.A1(_06318_),
    .A2(_05168_),
    .B1(_05388_),
    .B2(_05610_),
    .X(_07071_));
 sky130_fd_sc_hd__and4_2 _21390_ (.A(_06425_),
    .B(_11922_),
    .C(_06426_),
    .D(_11919_),
    .X(_07072_));
 sky130_fd_sc_hd__or2_2 _21391_ (.A(_07071_),
    .B(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__a2bb2o_2 _21392_ (.A1_N(_07070_),
    .A2_N(_07073_),
    .B1(_07070_),
    .B2(_07073_),
    .X(_07074_));
 sky130_fd_sc_hd__a2bb2o_2 _21393_ (.A1_N(_07069_),
    .A2_N(_07074_),
    .B1(_07069_),
    .B2(_07074_),
    .X(_07075_));
 sky130_fd_sc_hd__a2bb2o_2 _21394_ (.A1_N(_07068_),
    .A2_N(_07075_),
    .B1(_07068_),
    .B2(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__o22a_2 _21395_ (.A1(_06937_),
    .A2(_06942_),
    .B1(_06936_),
    .B2(_06943_),
    .X(_07077_));
 sky130_fd_sc_hd__a2bb2o_2 _21396_ (.A1_N(_07076_),
    .A2_N(_07077_),
    .B1(_07076_),
    .B2(_07077_),
    .X(_07078_));
 sky130_fd_sc_hd__a2bb2o_2 _21397_ (.A1_N(_07067_),
    .A2_N(_07078_),
    .B1(_07067_),
    .B2(_07078_),
    .X(_07079_));
 sky130_fd_sc_hd__a2bb2o_2 _21398_ (.A1_N(_07053_),
    .A2_N(_07079_),
    .B1(_07053_),
    .B2(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__a2bb2o_2 _21399_ (.A1_N(_07052_),
    .A2_N(_07080_),
    .B1(_07052_),
    .B2(_07080_),
    .X(_07081_));
 sky130_fd_sc_hd__o22a_2 _21400_ (.A1(_06960_),
    .A2(_06961_),
    .B1(_06955_),
    .B2(_06962_),
    .X(_07082_));
 sky130_fd_sc_hd__o22a_2 _21401_ (.A1(_06834_),
    .A2(_06978_),
    .B1(_06972_),
    .B2(_06979_),
    .X(_07083_));
 sky130_fd_sc_hd__or2_2 _21402_ (.A(_06451_),
    .B(_05937_),
    .X(_07084_));
 sky130_fd_sc_hd__o22a_2 _21403_ (.A1(_06572_),
    .A2(_05163_),
    .B1(_06573_),
    .B2(_05345_),
    .X(_07085_));
 sky130_fd_sc_hd__and4_2 _21404_ (.A(_06453_),
    .B(_05260_),
    .C(_06280_),
    .D(_11926_),
    .X(_07086_));
 sky130_fd_sc_hd__or2_2 _21405_ (.A(_07085_),
    .B(_07086_),
    .X(_07087_));
 sky130_fd_sc_hd__a2bb2o_2 _21406_ (.A1_N(_07084_),
    .A2_N(_07087_),
    .B1(_07084_),
    .B2(_07087_),
    .X(_07088_));
 sky130_fd_sc_hd__or2_2 _21407_ (.A(_06035_),
    .B(_05077_),
    .X(_07089_));
 sky130_fd_sc_hd__o22a_2 _21408_ (.A1(_06579_),
    .A2(_05575_),
    .B1(_06033_),
    .B2(_05273_),
    .X(_07090_));
 sky130_fd_sc_hd__and4_2 _21409_ (.A(_11585_),
    .B(_05577_),
    .C(_11589_),
    .D(_05176_),
    .X(_07091_));
 sky130_fd_sc_hd__or2_2 _21410_ (.A(_07090_),
    .B(_07091_),
    .X(_07092_));
 sky130_fd_sc_hd__a2bb2o_2 _21411_ (.A1_N(_07089_),
    .A2_N(_07092_),
    .B1(_07089_),
    .B2(_07092_),
    .X(_07093_));
 sky130_fd_sc_hd__o21ba_2 _21412_ (.A1(_06956_),
    .A2(_06959_),
    .B1_N(_06958_),
    .X(_07094_));
 sky130_fd_sc_hd__a2bb2o_2 _21413_ (.A1_N(_07093_),
    .A2_N(_07094_),
    .B1(_07093_),
    .B2(_07094_),
    .X(_07095_));
 sky130_fd_sc_hd__a2bb2o_2 _21414_ (.A1_N(_07088_),
    .A2_N(_07095_),
    .B1(_07088_),
    .B2(_07095_),
    .X(_07096_));
 sky130_fd_sc_hd__a2bb2o_2 _21415_ (.A1_N(_07083_),
    .A2_N(_07096_),
    .B1(_07083_),
    .B2(_07096_),
    .X(_07097_));
 sky130_fd_sc_hd__a2bb2o_2 _21416_ (.A1_N(_07082_),
    .A2_N(_07097_),
    .B1(_07082_),
    .B2(_07097_),
    .X(_07098_));
 sky130_vsdinv _21417_ (.A(\pcpi_mul.rs2[30] ),
    .Y(_07099_));
 sky130_fd_sc_hd__buf_1 _21418_ (.A(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__buf_1 _21419_ (.A(_07100_),
    .X(_07101_));
 sky130_fd_sc_hd__or2_2 _21420_ (.A(_07101_),
    .B(_04543_),
    .X(_07102_));
 sky130_fd_sc_hd__or2_2 _21421_ (.A(_06684_),
    .B(_04723_),
    .X(_07103_));
 sky130_fd_sc_hd__and4_2 _21422_ (.A(\pcpi_mul.rs2[29] ),
    .B(_11955_),
    .C(\pcpi_mul.rs2[28] ),
    .D(_05144_),
    .X(_07104_));
 sky130_fd_sc_hd__o22a_2 _21423_ (.A1(_06968_),
    .A2(_04751_),
    .B1(_06828_),
    .B2(_04779_),
    .X(_07105_));
 sky130_fd_sc_hd__or2_2 _21424_ (.A(_07104_),
    .B(_07105_),
    .X(_07106_));
 sky130_fd_sc_hd__a2bb2o_2 _21425_ (.A1_N(_07103_),
    .A2_N(_07106_),
    .B1(_07103_),
    .B2(_07106_),
    .X(_07107_));
 sky130_fd_sc_hd__or2_2 _21426_ (.A(_07102_),
    .B(_07107_),
    .X(_07108_));
 sky130_fd_sc_hd__a21bo_2 _21427_ (.A1(_07102_),
    .A2(_07107_),
    .B1_N(_07108_),
    .X(_07109_));
 sky130_fd_sc_hd__o21ba_2 _21428_ (.A1(_06973_),
    .A2(_06977_),
    .B1_N(_06976_),
    .X(_07110_));
 sky130_fd_sc_hd__o21ba_2 _21429_ (.A1(_06966_),
    .A2(_06970_),
    .B1_N(_06967_),
    .X(_07111_));
 sky130_fd_sc_hd__or2_2 _21430_ (.A(_06272_),
    .B(_05312_),
    .X(_07112_));
 sky130_fd_sc_hd__o22a_2 _21431_ (.A1(_06974_),
    .A2(_05227_),
    .B1(_06441_),
    .B2(_05314_),
    .X(_07113_));
 sky130_fd_sc_hd__and4_2 _21432_ (.A(_11574_),
    .B(_05316_),
    .C(_11579_),
    .D(_11942_),
    .X(_07114_));
 sky130_fd_sc_hd__or2_2 _21433_ (.A(_07113_),
    .B(_07114_),
    .X(_07115_));
 sky130_fd_sc_hd__a2bb2o_2 _21434_ (.A1_N(_07112_),
    .A2_N(_07115_),
    .B1(_07112_),
    .B2(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__a2bb2o_2 _21435_ (.A1_N(_07111_),
    .A2_N(_07116_),
    .B1(_07111_),
    .B2(_07116_),
    .X(_07117_));
 sky130_fd_sc_hd__a2bb2o_2 _21436_ (.A1_N(_07110_),
    .A2_N(_07117_),
    .B1(_07110_),
    .B2(_07117_),
    .X(_07118_));
 sky130_fd_sc_hd__or2_2 _21437_ (.A(_07109_),
    .B(_07118_),
    .X(_07119_));
 sky130_fd_sc_hd__a21bo_2 _21438_ (.A1(_07109_),
    .A2(_07118_),
    .B1_N(_07119_),
    .X(_07120_));
 sky130_fd_sc_hd__a2bb2o_2 _21439_ (.A1_N(_06981_),
    .A2_N(_07120_),
    .B1(_06981_),
    .B2(_07120_),
    .X(_07121_));
 sky130_fd_sc_hd__a2bb2o_2 _21440_ (.A1_N(_07098_),
    .A2_N(_07121_),
    .B1(_07098_),
    .B2(_07121_),
    .X(_07122_));
 sky130_fd_sc_hd__o22a_2 _21441_ (.A1(_06844_),
    .A2(_06982_),
    .B1(_06965_),
    .B2(_06983_),
    .X(_07123_));
 sky130_fd_sc_hd__a2bb2o_2 _21442_ (.A1_N(_07122_),
    .A2_N(_07123_),
    .B1(_07122_),
    .B2(_07123_),
    .X(_07124_));
 sky130_fd_sc_hd__a2bb2o_2 _21443_ (.A1_N(_07081_),
    .A2_N(_07124_),
    .B1(_07081_),
    .B2(_07124_),
    .X(_07125_));
 sky130_fd_sc_hd__o22a_2 _21444_ (.A1(_06984_),
    .A2(_06985_),
    .B1(_06949_),
    .B2(_06986_),
    .X(_07126_));
 sky130_fd_sc_hd__a2bb2o_2 _21445_ (.A1_N(_07125_),
    .A2_N(_07126_),
    .B1(_07125_),
    .B2(_07126_),
    .X(_07127_));
 sky130_fd_sc_hd__a2bb2o_2 _21446_ (.A1_N(_07051_),
    .A2_N(_07127_),
    .B1(_07051_),
    .B2(_07127_),
    .X(_07128_));
 sky130_fd_sc_hd__o22a_2 _21447_ (.A1(_06987_),
    .A2(_06988_),
    .B1(_06918_),
    .B2(_06989_),
    .X(_07129_));
 sky130_fd_sc_hd__a2bb2o_2 _21448_ (.A1_N(_07128_),
    .A2_N(_07129_),
    .B1(_07128_),
    .B2(_07129_),
    .X(_07130_));
 sky130_fd_sc_hd__a2bb2o_2 _21449_ (.A1_N(_07003_),
    .A2_N(_07130_),
    .B1(_07003_),
    .B2(_07130_),
    .X(_07131_));
 sky130_fd_sc_hd__o22a_2 _21450_ (.A1(_06990_),
    .A2(_06991_),
    .B1(_06872_),
    .B2(_06992_),
    .X(_07132_));
 sky130_fd_sc_hd__a2bb2o_2 _21451_ (.A1_N(_07131_),
    .A2_N(_07132_),
    .B1(_07131_),
    .B2(_07132_),
    .X(_07133_));
 sky130_fd_sc_hd__a2bb2o_2 _21452_ (.A1_N(_06871_),
    .A2_N(_07133_),
    .B1(_06871_),
    .B2(_07133_),
    .X(_07134_));
 sky130_fd_sc_hd__o22a_2 _21453_ (.A1(_06993_),
    .A2(_06994_),
    .B1(_06736_),
    .B2(_06995_),
    .X(_07135_));
 sky130_fd_sc_hd__or2_2 _21454_ (.A(_07134_),
    .B(_07135_),
    .X(_07136_));
 sky130_fd_sc_hd__a21bo_2 _21455_ (.A1(_07134_),
    .A2(_07135_),
    .B1_N(_07136_),
    .X(_07137_));
 sky130_fd_sc_hd__a22o_2 _21456_ (.A1(_06868_),
    .A2(_06996_),
    .B1(_06860_),
    .B2(_06997_),
    .X(_07138_));
 sky130_fd_sc_hd__o31a_2 _21457_ (.A1(_06861_),
    .A2(_06998_),
    .A3(_06866_),
    .B1(_07138_),
    .X(_07139_));
 sky130_fd_sc_hd__a2bb2oi_2 _21458_ (.A1_N(_07137_),
    .A2_N(_07139_),
    .B1(_07137_),
    .B2(_07139_),
    .Y(_02649_));
 sky130_fd_sc_hd__o22a_2 _21459_ (.A1(_07131_),
    .A2(_07132_),
    .B1(_06871_),
    .B2(_07133_),
    .X(_07140_));
 sky130_fd_sc_hd__o22a_2 _21460_ (.A1(_07005_),
    .A2(_07049_),
    .B1(_07004_),
    .B2(_07050_),
    .X(_07141_));
 sky130_fd_sc_hd__o22a_2 _21461_ (.A1(_07029_),
    .A2(_07030_),
    .B1(_07006_),
    .B2(_07031_),
    .X(_07142_));
 sky130_fd_sc_hd__or2_2 _21462_ (.A(_07141_),
    .B(_07142_),
    .X(_07143_));
 sky130_fd_sc_hd__a21bo_2 _21463_ (.A1(_07141_),
    .A2(_07142_),
    .B1_N(_07143_),
    .X(_07144_));
 sky130_fd_sc_hd__o22a_2 _21464_ (.A1(_07046_),
    .A2(_07047_),
    .B1(_07032_),
    .B2(_07048_),
    .X(_07145_));
 sky130_fd_sc_hd__o22a_2 _21465_ (.A1(_07053_),
    .A2(_07079_),
    .B1(_07052_),
    .B2(_07080_),
    .X(_07146_));
 sky130_fd_sc_hd__a21oi_2 _21466_ (.A1(_07014_),
    .A2(_07016_),
    .B1(_07013_),
    .Y(_07147_));
 sky130_fd_sc_hd__o22a_2 _21467_ (.A1(_05813_),
    .A2(_07010_),
    .B1(_05703_),
    .B2(_07024_),
    .X(_07148_));
 sky130_fd_sc_hd__and4_2 _21468_ (.A(_05706_),
    .B(_07012_),
    .C(_05707_),
    .D(_11878_),
    .X(_07149_));
 sky130_fd_sc_hd__nor2_2 _21469_ (.A(_07148_),
    .B(_07149_),
    .Y(_07150_));
 sky130_fd_sc_hd__buf_1 _21470_ (.A(_06750_),
    .X(_07151_));
 sky130_fd_sc_hd__nor2_2 _21471_ (.A(_05710_),
    .B(_07151_),
    .Y(_07152_));
 sky130_fd_sc_hd__a2bb2o_2 _21472_ (.A1_N(_07150_),
    .A2_N(_07152_),
    .B1(_07150_),
    .B2(_07152_),
    .X(_07153_));
 sky130_fd_sc_hd__o22a_2 _21473_ (.A1(_06368_),
    .A2(_06496_),
    .B1(_06369_),
    .B2(_06879_),
    .X(_07154_));
 sky130_fd_sc_hd__buf_1 _21474_ (.A(_11884_),
    .X(_07155_));
 sky130_fd_sc_hd__and4_2 _21475_ (.A(_11629_),
    .B(_11888_),
    .C(_11633_),
    .D(_07155_),
    .X(_07156_));
 sky130_fd_sc_hd__nor2_2 _21476_ (.A(_07154_),
    .B(_07156_),
    .Y(_07157_));
 sky130_vsdinv _21477_ (.A(\pcpi_mul.rs1[31] ),
    .Y(_07158_));
 sky130_fd_sc_hd__buf_1 _21478_ (.A(_07158_),
    .X(_07159_));
 sky130_fd_sc_hd__buf_1 _21479_ (.A(_07159_),
    .X(_07160_));
 sky130_fd_sc_hd__nor2_2 _21480_ (.A(_04538_),
    .B(_07160_),
    .Y(_07161_));
 sky130_fd_sc_hd__a2bb2o_2 _21481_ (.A1_N(_07157_),
    .A2_N(_07161_),
    .B1(_07157_),
    .B2(_07161_),
    .X(_07162_));
 sky130_fd_sc_hd__a21oi_2 _21482_ (.A1(_07020_),
    .A2(_07025_),
    .B1(_07019_),
    .Y(_07163_));
 sky130_fd_sc_hd__a2bb2o_2 _21483_ (.A1_N(_07162_),
    .A2_N(_07163_),
    .B1(_07162_),
    .B2(_07163_),
    .X(_07164_));
 sky130_fd_sc_hd__a2bb2o_2 _21484_ (.A1_N(_07153_),
    .A2_N(_07164_),
    .B1(_07153_),
    .B2(_07164_),
    .X(_07165_));
 sky130_fd_sc_hd__o22a_2 _21485_ (.A1(_07026_),
    .A2(_07027_),
    .B1(_07017_),
    .B2(_07028_),
    .X(_07166_));
 sky130_fd_sc_hd__a2bb2o_2 _21486_ (.A1_N(_07165_),
    .A2_N(_07166_),
    .B1(_07165_),
    .B2(_07166_),
    .X(_07167_));
 sky130_fd_sc_hd__a2bb2o_2 _21487_ (.A1_N(_07147_),
    .A2_N(_07167_),
    .B1(_07147_),
    .B2(_07167_),
    .X(_07168_));
 sky130_fd_sc_hd__o22a_2 _21488_ (.A1(_07036_),
    .A2(_07042_),
    .B1(_07035_),
    .B2(_07043_),
    .X(_07169_));
 sky130_fd_sc_hd__o22a_2 _21489_ (.A1(_07064_),
    .A2(_07065_),
    .B1(_07058_),
    .B2(_07066_),
    .X(_07170_));
 sky130_fd_sc_hd__a21oi_2 _21490_ (.A1(_07040_),
    .A2(_07041_),
    .B1(_07039_),
    .Y(_07171_));
 sky130_fd_sc_hd__o21ba_2 _21491_ (.A1(_07054_),
    .A2(_07057_),
    .B1_N(_07056_),
    .X(_07172_));
 sky130_fd_sc_hd__buf_1 _21492_ (.A(_06232_),
    .X(_07173_));
 sky130_fd_sc_hd__o22a_2 _21493_ (.A1(_06132_),
    .A2(_06111_),
    .B1(_06133_),
    .B2(_07173_),
    .X(_07174_));
 sky130_fd_sc_hd__buf_1 _21494_ (.A(\pcpi_mul.rs1[24] ),
    .X(_07175_));
 sky130_fd_sc_hd__and4_2 _21495_ (.A(_06136_),
    .B(_07038_),
    .C(_06137_),
    .D(_07175_),
    .X(_07176_));
 sky130_fd_sc_hd__nor2_2 _21496_ (.A(_07174_),
    .B(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__nor2_2 _21497_ (.A(_04830_),
    .B(_06377_),
    .Y(_07178_));
 sky130_fd_sc_hd__a2bb2o_2 _21498_ (.A1_N(_07177_),
    .A2_N(_07178_),
    .B1(_07177_),
    .B2(_07178_),
    .X(_07179_));
 sky130_fd_sc_hd__a2bb2o_2 _21499_ (.A1_N(_07172_),
    .A2_N(_07179_),
    .B1(_07172_),
    .B2(_07179_),
    .X(_07180_));
 sky130_fd_sc_hd__a2bb2o_2 _21500_ (.A1_N(_07171_),
    .A2_N(_07180_),
    .B1(_07171_),
    .B2(_07180_),
    .X(_07181_));
 sky130_fd_sc_hd__a2bb2o_2 _21501_ (.A1_N(_07170_),
    .A2_N(_07181_),
    .B1(_07170_),
    .B2(_07181_),
    .X(_07182_));
 sky130_fd_sc_hd__a2bb2o_2 _21502_ (.A1_N(_07169_),
    .A2_N(_07182_),
    .B1(_07169_),
    .B2(_07182_),
    .X(_07183_));
 sky130_fd_sc_hd__o22a_2 _21503_ (.A1(_07034_),
    .A2(_07044_),
    .B1(_07033_),
    .B2(_07045_),
    .X(_07184_));
 sky130_fd_sc_hd__a2bb2o_2 _21504_ (.A1_N(_07183_),
    .A2_N(_07184_),
    .B1(_07183_),
    .B2(_07184_),
    .X(_07185_));
 sky130_fd_sc_hd__a2bb2o_2 _21505_ (.A1_N(_07168_),
    .A2_N(_07185_),
    .B1(_07168_),
    .B2(_07185_),
    .X(_07186_));
 sky130_fd_sc_hd__a2bb2o_2 _21506_ (.A1_N(_07146_),
    .A2_N(_07186_),
    .B1(_07146_),
    .B2(_07186_),
    .X(_07187_));
 sky130_fd_sc_hd__a2bb2o_2 _21507_ (.A1_N(_07145_),
    .A2_N(_07187_),
    .B1(_07145_),
    .B2(_07187_),
    .X(_07188_));
 sky130_fd_sc_hd__o22a_2 _21508_ (.A1(_07076_),
    .A2(_07077_),
    .B1(_07067_),
    .B2(_07078_),
    .X(_07189_));
 sky130_fd_sc_hd__o22a_2 _21509_ (.A1(_07083_),
    .A2(_07096_),
    .B1(_07082_),
    .B2(_07097_),
    .X(_07190_));
 sky130_fd_sc_hd__or2_2 _21510_ (.A(_05665_),
    .B(_06502_),
    .X(_07191_));
 sky130_fd_sc_hd__o22a_2 _21511_ (.A1(_05779_),
    .A2(_06236_),
    .B1(_05667_),
    .B2(_05986_),
    .X(_07192_));
 sky130_fd_sc_hd__and4_2 _21512_ (.A(_05669_),
    .B(\pcpi_mul.rs1[20] ),
    .C(_05670_),
    .D(\pcpi_mul.rs1[21] ),
    .X(_07193_));
 sky130_fd_sc_hd__or2_2 _21513_ (.A(_07192_),
    .B(_07193_),
    .X(_07194_));
 sky130_fd_sc_hd__a2bb2o_2 _21514_ (.A1_N(_07191_),
    .A2_N(_07194_),
    .B1(_07191_),
    .B2(_07194_),
    .X(_07195_));
 sky130_fd_sc_hd__buf_1 _21515_ (.A(_05714_),
    .X(_07196_));
 sky130_fd_sc_hd__or2_2 _21516_ (.A(_05133_),
    .B(_07196_),
    .X(_07197_));
 sky130_fd_sc_hd__o22a_2 _21517_ (.A1(_05945_),
    .A2(_05509_),
    .B1(_06415_),
    .B2(_05606_),
    .X(_07198_));
 sky130_fd_sc_hd__and4_2 _21518_ (.A(_06928_),
    .B(_11912_),
    .C(_06929_),
    .D(_11910_),
    .X(_07199_));
 sky130_fd_sc_hd__or2_2 _21519_ (.A(_07198_),
    .B(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__a2bb2o_2 _21520_ (.A1_N(_07197_),
    .A2_N(_07200_),
    .B1(_07197_),
    .B2(_07200_),
    .X(_07201_));
 sky130_fd_sc_hd__o21ba_2 _21521_ (.A1(_07060_),
    .A2(_07063_),
    .B1_N(_07062_),
    .X(_07202_));
 sky130_fd_sc_hd__a2bb2o_2 _21522_ (.A1_N(_07201_),
    .A2_N(_07202_),
    .B1(_07201_),
    .B2(_07202_),
    .X(_07203_));
 sky130_fd_sc_hd__a2bb2o_2 _21523_ (.A1_N(_07195_),
    .A2_N(_07203_),
    .B1(_07195_),
    .B2(_07203_),
    .X(_07204_));
 sky130_fd_sc_hd__o21ba_2 _21524_ (.A1(_07070_),
    .A2(_07073_),
    .B1_N(_07072_),
    .X(_07205_));
 sky130_fd_sc_hd__o21ba_2 _21525_ (.A1(_07084_),
    .A2(_07087_),
    .B1_N(_07086_),
    .X(_07206_));
 sky130_fd_sc_hd__or2_2 _21526_ (.A(_05393_),
    .B(_05429_),
    .X(_07207_));
 sky130_fd_sc_hd__o22a_2 _21527_ (.A1(_06318_),
    .A2(_05255_),
    .B1(_05388_),
    .B2(_06014_),
    .X(_07208_));
 sky130_fd_sc_hd__and4_2 _21528_ (.A(_11602_),
    .B(_11919_),
    .C(_11605_),
    .D(_11916_),
    .X(_07209_));
 sky130_fd_sc_hd__or2_2 _21529_ (.A(_07208_),
    .B(_07209_),
    .X(_07210_));
 sky130_fd_sc_hd__a2bb2o_2 _21530_ (.A1_N(_07207_),
    .A2_N(_07210_),
    .B1(_07207_),
    .B2(_07210_),
    .X(_07211_));
 sky130_fd_sc_hd__a2bb2o_2 _21531_ (.A1_N(_07206_),
    .A2_N(_07211_),
    .B1(_07206_),
    .B2(_07211_),
    .X(_07212_));
 sky130_fd_sc_hd__a2bb2o_2 _21532_ (.A1_N(_07205_),
    .A2_N(_07212_),
    .B1(_07205_),
    .B2(_07212_),
    .X(_07213_));
 sky130_fd_sc_hd__o22a_2 _21533_ (.A1(_07069_),
    .A2(_07074_),
    .B1(_07068_),
    .B2(_07075_),
    .X(_07214_));
 sky130_fd_sc_hd__a2bb2o_2 _21534_ (.A1_N(_07213_),
    .A2_N(_07214_),
    .B1(_07213_),
    .B2(_07214_),
    .X(_07215_));
 sky130_fd_sc_hd__a2bb2o_2 _21535_ (.A1_N(_07204_),
    .A2_N(_07215_),
    .B1(_07204_),
    .B2(_07215_),
    .X(_07216_));
 sky130_fd_sc_hd__a2bb2o_2 _21536_ (.A1_N(_07190_),
    .A2_N(_07216_),
    .B1(_07190_),
    .B2(_07216_),
    .X(_07217_));
 sky130_fd_sc_hd__a2bb2o_2 _21537_ (.A1_N(_07189_),
    .A2_N(_07217_),
    .B1(_07189_),
    .B2(_07217_),
    .X(_07218_));
 sky130_fd_sc_hd__o22a_2 _21538_ (.A1(_07093_),
    .A2(_07094_),
    .B1(_07088_),
    .B2(_07095_),
    .X(_07219_));
 sky130_fd_sc_hd__o22a_2 _21539_ (.A1(_07111_),
    .A2(_07116_),
    .B1(_07110_),
    .B2(_07117_),
    .X(_07220_));
 sky130_fd_sc_hd__or2_2 _21540_ (.A(_06451_),
    .B(_05736_),
    .X(_07221_));
 sky130_fd_sc_hd__o22a_2 _21541_ (.A1(_06572_),
    .A2(_05345_),
    .B1(_06573_),
    .B2(_05431_),
    .X(_07222_));
 sky130_fd_sc_hd__and4_2 _21542_ (.A(_06453_),
    .B(_05433_),
    .C(_06280_),
    .D(_11924_),
    .X(_07223_));
 sky130_fd_sc_hd__or2_2 _21543_ (.A(_07222_),
    .B(_07223_),
    .X(_07224_));
 sky130_fd_sc_hd__a2bb2o_2 _21544_ (.A1_N(_07221_),
    .A2_N(_07224_),
    .B1(_07221_),
    .B2(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__or2_2 _21545_ (.A(_05926_),
    .B(_05164_),
    .X(_07226_));
 sky130_fd_sc_hd__o22a_2 _21546_ (.A1(_06818_),
    .A2(_05172_),
    .B1(_06033_),
    .B2(_06429_),
    .X(_07227_));
 sky130_fd_sc_hd__and4_2 _21547_ (.A(_11585_),
    .B(_05176_),
    .C(_11589_),
    .D(_05781_),
    .X(_07228_));
 sky130_fd_sc_hd__or2_2 _21548_ (.A(_07227_),
    .B(_07228_),
    .X(_07229_));
 sky130_fd_sc_hd__a2bb2o_2 _21549_ (.A1_N(_07226_),
    .A2_N(_07229_),
    .B1(_07226_),
    .B2(_07229_),
    .X(_07230_));
 sky130_fd_sc_hd__o21ba_2 _21550_ (.A1(_07089_),
    .A2(_07092_),
    .B1_N(_07091_),
    .X(_07231_));
 sky130_fd_sc_hd__a2bb2o_2 _21551_ (.A1_N(_07230_),
    .A2_N(_07231_),
    .B1(_07230_),
    .B2(_07231_),
    .X(_07232_));
 sky130_fd_sc_hd__a2bb2o_2 _21552_ (.A1_N(_07225_),
    .A2_N(_07232_),
    .B1(_07225_),
    .B2(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__a2bb2o_2 _21553_ (.A1_N(_07220_),
    .A2_N(_07233_),
    .B1(_07220_),
    .B2(_07233_),
    .X(_07234_));
 sky130_fd_sc_hd__a2bb2o_2 _21554_ (.A1_N(_07219_),
    .A2_N(_07234_),
    .B1(_07219_),
    .B2(_07234_),
    .X(_07235_));
 sky130_fd_sc_hd__o21ba_2 _21555_ (.A1(_07112_),
    .A2(_07115_),
    .B1_N(_07114_),
    .X(_07236_));
 sky130_fd_sc_hd__o21ba_2 _21556_ (.A1(_07103_),
    .A2(_07106_),
    .B1_N(_07104_),
    .X(_07237_));
 sky130_fd_sc_hd__or2_2 _21557_ (.A(_06272_),
    .B(_05191_),
    .X(_07238_));
 sky130_fd_sc_hd__o22a_2 _21558_ (.A1(_06974_),
    .A2(_05225_),
    .B1(_06441_),
    .B2(_06277_),
    .X(_07239_));
 sky130_fd_sc_hd__buf_1 _21559_ (.A(_11574_),
    .X(_07240_));
 sky130_fd_sc_hd__and4_2 _21560_ (.A(_07240_),
    .B(_11943_),
    .C(_11580_),
    .D(_11940_),
    .X(_07241_));
 sky130_fd_sc_hd__or2_2 _21561_ (.A(_07239_),
    .B(_07241_),
    .X(_07242_));
 sky130_fd_sc_hd__a2bb2o_2 _21562_ (.A1_N(_07238_),
    .A2_N(_07242_),
    .B1(_07238_),
    .B2(_07242_),
    .X(_07243_));
 sky130_fd_sc_hd__a2bb2o_2 _21563_ (.A1_N(_07237_),
    .A2_N(_07243_),
    .B1(_07237_),
    .B2(_07243_),
    .X(_07244_));
 sky130_fd_sc_hd__a2bb2o_2 _21564_ (.A1_N(_07236_),
    .A2_N(_07244_),
    .B1(_07236_),
    .B2(_07244_),
    .X(_07245_));
 sky130_vsdinv _21565_ (.A(\pcpi_mul.rs2[31] ),
    .Y(_07246_));
 sky130_fd_sc_hd__buf_1 _21566_ (.A(_07246_),
    .X(_07247_));
 sky130_fd_sc_hd__o22a_2 _21567_ (.A1(_07247_),
    .A2(_04542_),
    .B1(_07100_),
    .B2(_04703_),
    .X(_07248_));
 sky130_fd_sc_hd__or4_2 _21568_ (.A(_07247_),
    .B(_04542_),
    .C(_07099_),
    .D(_04688_),
    .X(_07249_));
 sky130_fd_sc_hd__or2b_2 _21569_ (.A(_07248_),
    .B_N(_07249_),
    .X(_07250_));
 sky130_fd_sc_hd__or2_2 _21570_ (.A(_06684_),
    .B(_05403_),
    .X(_07251_));
 sky130_fd_sc_hd__and4_2 _21571_ (.A(_11566_),
    .B(_11952_),
    .C(_11570_),
    .D(_05145_),
    .X(_07252_));
 sky130_fd_sc_hd__o22a_2 _21572_ (.A1(_06968_),
    .A2(_05061_),
    .B1(_06828_),
    .B2(_05141_),
    .X(_07253_));
 sky130_fd_sc_hd__or2_2 _21573_ (.A(_07252_),
    .B(_07253_),
    .X(_07254_));
 sky130_fd_sc_hd__a2bb2o_2 _21574_ (.A1_N(_07251_),
    .A2_N(_07254_),
    .B1(_07251_),
    .B2(_07254_),
    .X(_07255_));
 sky130_fd_sc_hd__or2_2 _21575_ (.A(_07250_),
    .B(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__a21bo_2 _21576_ (.A1(_07250_),
    .A2(_07255_),
    .B1_N(_07256_),
    .X(_07257_));
 sky130_fd_sc_hd__a2bb2o_2 _21577_ (.A1_N(_07108_),
    .A2_N(_07257_),
    .B1(_07108_),
    .B2(_07257_),
    .X(_07258_));
 sky130_fd_sc_hd__a2bb2o_2 _21578_ (.A1_N(_07245_),
    .A2_N(_07258_),
    .B1(_07245_),
    .B2(_07258_),
    .X(_07259_));
 sky130_fd_sc_hd__a2bb2o_2 _21579_ (.A1_N(_07119_),
    .A2_N(_07259_),
    .B1(_07119_),
    .B2(_07259_),
    .X(_07260_));
 sky130_fd_sc_hd__a2bb2o_2 _21580_ (.A1_N(_07235_),
    .A2_N(_07260_),
    .B1(_07235_),
    .B2(_07260_),
    .X(_07261_));
 sky130_fd_sc_hd__o22a_2 _21581_ (.A1(_06981_),
    .A2(_07120_),
    .B1(_07098_),
    .B2(_07121_),
    .X(_07262_));
 sky130_fd_sc_hd__a2bb2o_2 _21582_ (.A1_N(_07261_),
    .A2_N(_07262_),
    .B1(_07261_),
    .B2(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__a2bb2o_2 _21583_ (.A1_N(_07218_),
    .A2_N(_07263_),
    .B1(_07218_),
    .B2(_07263_),
    .X(_07264_));
 sky130_fd_sc_hd__o22a_2 _21584_ (.A1(_07122_),
    .A2(_07123_),
    .B1(_07081_),
    .B2(_07124_),
    .X(_07265_));
 sky130_fd_sc_hd__a2bb2o_2 _21585_ (.A1_N(_07264_),
    .A2_N(_07265_),
    .B1(_07264_),
    .B2(_07265_),
    .X(_07266_));
 sky130_fd_sc_hd__a2bb2o_2 _21586_ (.A1_N(_07188_),
    .A2_N(_07266_),
    .B1(_07188_),
    .B2(_07266_),
    .X(_07267_));
 sky130_fd_sc_hd__o22a_2 _21587_ (.A1(_07125_),
    .A2(_07126_),
    .B1(_07051_),
    .B2(_07127_),
    .X(_07268_));
 sky130_fd_sc_hd__a2bb2o_2 _21588_ (.A1_N(_07267_),
    .A2_N(_07268_),
    .B1(_07267_),
    .B2(_07268_),
    .X(_07269_));
 sky130_fd_sc_hd__a2bb2o_2 _21589_ (.A1_N(_07144_),
    .A2_N(_07269_),
    .B1(_07144_),
    .B2(_07269_),
    .X(_07270_));
 sky130_fd_sc_hd__o22a_2 _21590_ (.A1(_07128_),
    .A2(_07129_),
    .B1(_07003_),
    .B2(_07130_),
    .X(_07271_));
 sky130_fd_sc_hd__a2bb2o_2 _21591_ (.A1_N(_07270_),
    .A2_N(_07271_),
    .B1(_07270_),
    .B2(_07271_),
    .X(_07272_));
 sky130_fd_sc_hd__a2bb2o_2 _21592_ (.A1_N(_07002_),
    .A2_N(_07272_),
    .B1(_07002_),
    .B2(_07272_),
    .X(_07273_));
 sky130_fd_sc_hd__and2_2 _21593_ (.A(_07140_),
    .B(_07273_),
    .X(_07274_));
 sky130_fd_sc_hd__or2_2 _21594_ (.A(_07140_),
    .B(_07273_),
    .X(_07275_));
 sky130_fd_sc_hd__or2b_2 _21595_ (.A(_07274_),
    .B_N(_07275_),
    .X(_07276_));
 sky130_fd_sc_hd__o21ai_2 _21596_ (.A1(_07137_),
    .A2(_07139_),
    .B1(_07136_),
    .Y(_07277_));
 sky130_fd_sc_hd__a2bb2o_2 _21597_ (.A1_N(_07276_),
    .A2_N(_07277_),
    .B1(_07276_),
    .B2(_07277_),
    .X(_02650_));
 sky130_fd_sc_hd__o22a_2 _21598_ (.A1(_07146_),
    .A2(_07186_),
    .B1(_07145_),
    .B2(_07187_),
    .X(_07278_));
 sky130_fd_sc_hd__o22a_2 _21599_ (.A1(_07165_),
    .A2(_07166_),
    .B1(_07147_),
    .B2(_07167_),
    .X(_07279_));
 sky130_fd_sc_hd__a2bb2o_2 _21600_ (.A1_N(_07278_),
    .A2_N(_07279_),
    .B1(_07278_),
    .B2(_07279_),
    .X(_07280_));
 sky130_fd_sc_hd__a2bb2o_2 _21601_ (.A1_N(_10600_),
    .A2_N(_07280_),
    .B1(_10600_),
    .B2(_07280_),
    .X(_07281_));
 sky130_fd_sc_hd__o22a_2 _21602_ (.A1(_07183_),
    .A2(_07184_),
    .B1(_07168_),
    .B2(_07185_),
    .X(_07282_));
 sky130_fd_sc_hd__o22a_2 _21603_ (.A1(_07190_),
    .A2(_07216_),
    .B1(_07189_),
    .B2(_07217_),
    .X(_07283_));
 sky130_fd_sc_hd__a21oi_2 _21604_ (.A1(_07150_),
    .A2(_07152_),
    .B1(_07149_),
    .Y(_07284_));
 sky130_fd_sc_hd__buf_1 _21605_ (.A(_07023_),
    .X(_07285_));
 sky130_fd_sc_hd__o22a_2 _21606_ (.A1(_05813_),
    .A2(_07285_),
    .B1(_05703_),
    .B2(_07160_),
    .X(_07286_));
 sky130_fd_sc_hd__and4_2 _21607_ (.A(_05706_),
    .B(_11877_),
    .C(_05707_),
    .D(_11874_),
    .X(_07287_));
 sky130_fd_sc_hd__nor2_2 _21608_ (.A(_07286_),
    .B(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__buf_1 _21609_ (.A(_06891_),
    .X(_07289_));
 sky130_fd_sc_hd__nor2_2 _21610_ (.A(_05710_),
    .B(_07289_),
    .Y(_07290_));
 sky130_fd_sc_hd__a2bb2o_2 _21611_ (.A1_N(_07288_),
    .A2_N(_07290_),
    .B1(_07288_),
    .B2(_07290_),
    .X(_07291_));
 sky130_fd_sc_hd__o22a_2 _21612_ (.A1(_06368_),
    .A2(_06624_),
    .B1(_06369_),
    .B2(_06750_),
    .X(_07292_));
 sky130_fd_sc_hd__and4_2 _21613_ (.A(_11629_),
    .B(_07155_),
    .C(_11633_),
    .D(_11882_),
    .X(_07293_));
 sky130_fd_sc_hd__nor2_2 _21614_ (.A(_07292_),
    .B(_07293_),
    .Y(_07294_));
 sky130_fd_sc_hd__or2_2 _21615_ (.A(_10585_),
    .B(_04536_),
    .X(_07295_));
 sky130_vsdinv _21616_ (.A(_07295_),
    .Y(_07296_));
 sky130_fd_sc_hd__buf_1 _21617_ (.A(_07296_),
    .X(_07297_));
 sky130_fd_sc_hd__a2bb2o_2 _21618_ (.A1_N(_07294_),
    .A2_N(_07297_),
    .B1(_07294_),
    .B2(_07297_),
    .X(_07298_));
 sky130_fd_sc_hd__a21oi_2 _21619_ (.A1(_07157_),
    .A2(_07161_),
    .B1(_07156_),
    .Y(_07299_));
 sky130_fd_sc_hd__a2bb2o_2 _21620_ (.A1_N(_07298_),
    .A2_N(_07299_),
    .B1(_07298_),
    .B2(_07299_),
    .X(_07300_));
 sky130_fd_sc_hd__a2bb2o_2 _21621_ (.A1_N(_07291_),
    .A2_N(_07300_),
    .B1(_07291_),
    .B2(_07300_),
    .X(_07301_));
 sky130_fd_sc_hd__o22a_2 _21622_ (.A1(_07162_),
    .A2(_07163_),
    .B1(_07153_),
    .B2(_07164_),
    .X(_07302_));
 sky130_fd_sc_hd__a2bb2o_2 _21623_ (.A1_N(_07301_),
    .A2_N(_07302_),
    .B1(_07301_),
    .B2(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__a2bb2o_2 _21624_ (.A1_N(_07284_),
    .A2_N(_07303_),
    .B1(_07284_),
    .B2(_07303_),
    .X(_07304_));
 sky130_fd_sc_hd__o22a_2 _21625_ (.A1(_07172_),
    .A2(_07179_),
    .B1(_07171_),
    .B2(_07180_),
    .X(_07305_));
 sky130_fd_sc_hd__o22a_2 _21626_ (.A1(_07201_),
    .A2(_07202_),
    .B1(_07195_),
    .B2(_07203_),
    .X(_07306_));
 sky130_fd_sc_hd__a21oi_2 _21627_ (.A1(_07177_),
    .A2(_07178_),
    .B1(_07176_),
    .Y(_07307_));
 sky130_fd_sc_hd__o21ba_2 _21628_ (.A1(_07191_),
    .A2(_07194_),
    .B1_N(_07193_),
    .X(_07308_));
 sky130_fd_sc_hd__o22a_2 _21629_ (.A1(_06132_),
    .A2(_07173_),
    .B1(_06133_),
    .B2(_06376_),
    .X(_07309_));
 sky130_fd_sc_hd__and4_2 _21630_ (.A(_06136_),
    .B(_07175_),
    .C(_06137_),
    .D(_11892_),
    .X(_07310_));
 sky130_fd_sc_hd__nor2_2 _21631_ (.A(_07309_),
    .B(_07310_),
    .Y(_07311_));
 sky130_fd_sc_hd__nor2_2 _21632_ (.A(_04830_),
    .B(_06743_),
    .Y(_07312_));
 sky130_fd_sc_hd__a2bb2o_2 _21633_ (.A1_N(_07311_),
    .A2_N(_07312_),
    .B1(_07311_),
    .B2(_07312_),
    .X(_07313_));
 sky130_fd_sc_hd__a2bb2o_2 _21634_ (.A1_N(_07308_),
    .A2_N(_07313_),
    .B1(_07308_),
    .B2(_07313_),
    .X(_07314_));
 sky130_fd_sc_hd__a2bb2o_2 _21635_ (.A1_N(_07307_),
    .A2_N(_07314_),
    .B1(_07307_),
    .B2(_07314_),
    .X(_07315_));
 sky130_fd_sc_hd__a2bb2o_2 _21636_ (.A1_N(_07306_),
    .A2_N(_07315_),
    .B1(_07306_),
    .B2(_07315_),
    .X(_07316_));
 sky130_fd_sc_hd__a2bb2o_2 _21637_ (.A1_N(_07305_),
    .A2_N(_07316_),
    .B1(_07305_),
    .B2(_07316_),
    .X(_07317_));
 sky130_fd_sc_hd__o22a_2 _21638_ (.A1(_07170_),
    .A2(_07181_),
    .B1(_07169_),
    .B2(_07182_),
    .X(_07318_));
 sky130_fd_sc_hd__a2bb2o_2 _21639_ (.A1_N(_07317_),
    .A2_N(_07318_),
    .B1(_07317_),
    .B2(_07318_),
    .X(_07319_));
 sky130_fd_sc_hd__a2bb2o_2 _21640_ (.A1_N(_07304_),
    .A2_N(_07319_),
    .B1(_07304_),
    .B2(_07319_),
    .X(_07320_));
 sky130_fd_sc_hd__a2bb2o_2 _21641_ (.A1_N(_07283_),
    .A2_N(_07320_),
    .B1(_07283_),
    .B2(_07320_),
    .X(_07321_));
 sky130_fd_sc_hd__a2bb2o_2 _21642_ (.A1_N(_07282_),
    .A2_N(_07321_),
    .B1(_07282_),
    .B2(_07321_),
    .X(_07322_));
 sky130_fd_sc_hd__o22a_2 _21643_ (.A1(_07213_),
    .A2(_07214_),
    .B1(_07204_),
    .B2(_07215_),
    .X(_07323_));
 sky130_fd_sc_hd__o22a_2 _21644_ (.A1(_07220_),
    .A2(_07233_),
    .B1(_07219_),
    .B2(_07234_),
    .X(_07324_));
 sky130_fd_sc_hd__or2_2 _21645_ (.A(_05665_),
    .B(_06359_),
    .X(_07325_));
 sky130_fd_sc_hd__o22a_2 _21646_ (.A1(_06299_),
    .A2(_05986_),
    .B1(_06300_),
    .B2(_05995_),
    .X(_07326_));
 sky130_fd_sc_hd__and4_2 _21647_ (.A(_06171_),
    .B(_06371_),
    .C(_06172_),
    .D(\pcpi_mul.rs1[22] ),
    .X(_07327_));
 sky130_fd_sc_hd__or2_2 _21648_ (.A(_07326_),
    .B(_07327_),
    .X(_07328_));
 sky130_fd_sc_hd__a2bb2o_2 _21649_ (.A1_N(_07325_),
    .A2_N(_07328_),
    .B1(_07325_),
    .B2(_07328_),
    .X(_07329_));
 sky130_fd_sc_hd__or2_2 _21650_ (.A(_06176_),
    .B(_05884_),
    .X(_07330_));
 sky130_fd_sc_hd__o22a_2 _21651_ (.A1(_06307_),
    .A2(_05606_),
    .B1(_06179_),
    .B2(_05814_),
    .X(_07331_));
 sky130_fd_sc_hd__and4_2 _21652_ (.A(_06928_),
    .B(_11910_),
    .C(_06929_),
    .D(_06517_),
    .X(_07332_));
 sky130_fd_sc_hd__or2_2 _21653_ (.A(_07331_),
    .B(_07332_),
    .X(_07333_));
 sky130_fd_sc_hd__a2bb2o_2 _21654_ (.A1_N(_07330_),
    .A2_N(_07333_),
    .B1(_07330_),
    .B2(_07333_),
    .X(_07334_));
 sky130_fd_sc_hd__o21ba_2 _21655_ (.A1(_07197_),
    .A2(_07200_),
    .B1_N(_07199_),
    .X(_07335_));
 sky130_fd_sc_hd__a2bb2o_2 _21656_ (.A1_N(_07334_),
    .A2_N(_07335_),
    .B1(_07334_),
    .B2(_07335_),
    .X(_07336_));
 sky130_fd_sc_hd__a2bb2o_2 _21657_ (.A1_N(_07329_),
    .A2_N(_07336_),
    .B1(_07329_),
    .B2(_07336_),
    .X(_07337_));
 sky130_fd_sc_hd__o21ba_2 _21658_ (.A1(_07207_),
    .A2(_07210_),
    .B1_N(_07209_),
    .X(_07338_));
 sky130_fd_sc_hd__o21ba_2 _21659_ (.A1(_07221_),
    .A2(_07224_),
    .B1_N(_07223_),
    .X(_07339_));
 sky130_fd_sc_hd__buf_1 _21660_ (.A(_06318_),
    .X(_07340_));
 sky130_fd_sc_hd__o22a_2 _21661_ (.A1(_07340_),
    .A2(_05420_),
    .B1(_05392_),
    .B2(_06134_),
    .X(_07341_));
 sky130_fd_sc_hd__buf_1 _21662_ (.A(_11602_),
    .X(_07342_));
 sky130_fd_sc_hd__buf_1 _21663_ (.A(_11605_),
    .X(_07343_));
 sky130_fd_sc_hd__and4_2 _21664_ (.A(_07342_),
    .B(_05830_),
    .C(_07343_),
    .D(_05831_),
    .X(_07344_));
 sky130_fd_sc_hd__nor2_2 _21665_ (.A(_07341_),
    .B(_07344_),
    .Y(_07345_));
 sky130_fd_sc_hd__buf_1 _21666_ (.A(_05308_),
    .X(_07346_));
 sky130_fd_sc_hd__nor2_2 _21667_ (.A(_07346_),
    .B(_05599_),
    .Y(_07347_));
 sky130_fd_sc_hd__a2bb2o_2 _21668_ (.A1_N(_07345_),
    .A2_N(_07347_),
    .B1(_07345_),
    .B2(_07347_),
    .X(_07348_));
 sky130_fd_sc_hd__a2bb2o_2 _21669_ (.A1_N(_07339_),
    .A2_N(_07348_),
    .B1(_07339_),
    .B2(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__a2bb2o_2 _21670_ (.A1_N(_07338_),
    .A2_N(_07349_),
    .B1(_07338_),
    .B2(_07349_),
    .X(_07350_));
 sky130_fd_sc_hd__o22a_2 _21671_ (.A1(_07206_),
    .A2(_07211_),
    .B1(_07205_),
    .B2(_07212_),
    .X(_07351_));
 sky130_fd_sc_hd__a2bb2o_2 _21672_ (.A1_N(_07350_),
    .A2_N(_07351_),
    .B1(_07350_),
    .B2(_07351_),
    .X(_07352_));
 sky130_fd_sc_hd__a2bb2o_2 _21673_ (.A1_N(_07337_),
    .A2_N(_07352_),
    .B1(_07337_),
    .B2(_07352_),
    .X(_07353_));
 sky130_fd_sc_hd__a2bb2o_2 _21674_ (.A1_N(_07324_),
    .A2_N(_07353_),
    .B1(_07324_),
    .B2(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__a2bb2o_2 _21675_ (.A1_N(_07323_),
    .A2_N(_07354_),
    .B1(_07323_),
    .B2(_07354_),
    .X(_07355_));
 sky130_fd_sc_hd__o22a_2 _21676_ (.A1(_07230_),
    .A2(_07231_),
    .B1(_07225_),
    .B2(_07232_),
    .X(_07356_));
 sky130_fd_sc_hd__o22a_2 _21677_ (.A1(_07237_),
    .A2(_07243_),
    .B1(_07236_),
    .B2(_07244_),
    .X(_07357_));
 sky130_fd_sc_hd__or2_2 _21678_ (.A(_06700_),
    .B(_05845_),
    .X(_07358_));
 sky130_fd_sc_hd__buf_1 _21679_ (.A(_06039_),
    .X(_07359_));
 sky130_fd_sc_hd__o22a_2 _21680_ (.A1(_07359_),
    .A2(_05157_),
    .B1(_05662_),
    .B2(_05246_),
    .X(_07360_));
 sky130_fd_sc_hd__and4_2 _21681_ (.A(_06703_),
    .B(_05745_),
    .C(_06570_),
    .D(_05848_),
    .X(_07361_));
 sky130_fd_sc_hd__or2_2 _21682_ (.A(_07360_),
    .B(_07361_),
    .X(_07362_));
 sky130_fd_sc_hd__a2bb2o_2 _21683_ (.A1_N(_07358_),
    .A2_N(_07362_),
    .B1(_07358_),
    .B2(_07362_),
    .X(_07363_));
 sky130_fd_sc_hd__or2_2 _21684_ (.A(_05926_),
    .B(_05155_),
    .X(_07364_));
 sky130_fd_sc_hd__o22a_2 _21685_ (.A1(_06818_),
    .A2(_06429_),
    .B1(_06030_),
    .B2(_06180_),
    .X(_07365_));
 sky130_fd_sc_hd__and4_2 _21686_ (.A(_11585_),
    .B(_11931_),
    .C(_11589_),
    .D(_06184_),
    .X(_07366_));
 sky130_fd_sc_hd__or2_2 _21687_ (.A(_07365_),
    .B(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__a2bb2o_2 _21688_ (.A1_N(_07364_),
    .A2_N(_07367_),
    .B1(_07364_),
    .B2(_07367_),
    .X(_07368_));
 sky130_fd_sc_hd__o21ba_2 _21689_ (.A1(_07226_),
    .A2(_07229_),
    .B1_N(_07228_),
    .X(_07369_));
 sky130_fd_sc_hd__a2bb2o_2 _21690_ (.A1_N(_07368_),
    .A2_N(_07369_),
    .B1(_07368_),
    .B2(_07369_),
    .X(_07370_));
 sky130_fd_sc_hd__a2bb2o_2 _21691_ (.A1_N(_07363_),
    .A2_N(_07370_),
    .B1(_07363_),
    .B2(_07370_),
    .X(_07371_));
 sky130_fd_sc_hd__a2bb2o_2 _21692_ (.A1_N(_07357_),
    .A2_N(_07371_),
    .B1(_07357_),
    .B2(_07371_),
    .X(_07372_));
 sky130_fd_sc_hd__a2bb2o_2 _21693_ (.A1_N(_07356_),
    .A2_N(_07372_),
    .B1(_07356_),
    .B2(_07372_),
    .X(_07373_));
 sky130_fd_sc_hd__o21ba_2 _21694_ (.A1(_07238_),
    .A2(_07242_),
    .B1_N(_07241_),
    .X(_07374_));
 sky130_fd_sc_hd__o21ba_2 _21695_ (.A1(_07251_),
    .A2(_07254_),
    .B1_N(_07252_),
    .X(_07375_));
 sky130_fd_sc_hd__buf_1 _21696_ (.A(_06272_),
    .X(_07376_));
 sky130_fd_sc_hd__or2_2 _21697_ (.A(_07376_),
    .B(_06568_),
    .X(_07377_));
 sky130_fd_sc_hd__buf_1 _21698_ (.A(_06974_),
    .X(_07378_));
 sky130_fd_sc_hd__buf_1 _21699_ (.A(_06441_),
    .X(_07379_));
 sky130_fd_sc_hd__o22a_2 _21700_ (.A1(_07378_),
    .A2(_05312_),
    .B1(_07379_),
    .B2(_05396_),
    .X(_07380_));
 sky130_fd_sc_hd__and4_2 _21701_ (.A(_07240_),
    .B(_11940_),
    .C(_11580_),
    .D(_11937_),
    .X(_07381_));
 sky130_fd_sc_hd__or2_2 _21702_ (.A(_07380_),
    .B(_07381_),
    .X(_07382_));
 sky130_fd_sc_hd__a2bb2o_2 _21703_ (.A1_N(_07377_),
    .A2_N(_07382_),
    .B1(_07377_),
    .B2(_07382_),
    .X(_07383_));
 sky130_fd_sc_hd__a2bb2o_2 _21704_ (.A1_N(_07375_),
    .A2_N(_07383_),
    .B1(_07375_),
    .B2(_07383_),
    .X(_07384_));
 sky130_fd_sc_hd__a2bb2o_2 _21705_ (.A1_N(_07374_),
    .A2_N(_07384_),
    .B1(_07374_),
    .B2(_07384_),
    .X(_07385_));
 sky130_fd_sc_hd__or2_2 _21706_ (.A(_06685_),
    .B(_06151_),
    .X(_07386_));
 sky130_fd_sc_hd__buf_1 _21707_ (.A(_06968_),
    .X(_07387_));
 sky130_fd_sc_hd__o22a_2 _21708_ (.A1(_07387_),
    .A2(_04723_),
    .B1(_06829_),
    .B2(_05403_),
    .X(_07388_));
 sky130_fd_sc_hd__and4_2 _21709_ (.A(_11566_),
    .B(_11949_),
    .C(_11570_),
    .D(_11946_),
    .X(_07389_));
 sky130_fd_sc_hd__or2_2 _21710_ (.A(_07388_),
    .B(_07389_),
    .X(_07390_));
 sky130_fd_sc_hd__a2bb2o_2 _21711_ (.A1_N(_07386_),
    .A2_N(_07390_),
    .B1(_07386_),
    .B2(_07390_),
    .X(_07391_));
 sky130_fd_sc_hd__or2_2 _21712_ (.A(_07100_),
    .B(_04702_),
    .X(_07392_));
 sky130_fd_sc_hd__buf_1 _21713_ (.A(\pcpi_mul.rs2[32] ),
    .X(_07393_));
 sky130_fd_sc_hd__and4_2 _21714_ (.A(_11559_),
    .B(_11955_),
    .C(_07393_),
    .D(_04710_),
    .X(_07394_));
 sky130_fd_sc_hd__o22a_2 _21715_ (.A1(_07246_),
    .A2(_04709_),
    .B1(_10596_),
    .B2(_11957_),
    .X(_07395_));
 sky130_fd_sc_hd__or2_2 _21716_ (.A(_07394_),
    .B(_07395_),
    .X(_07396_));
 sky130_fd_sc_hd__a2bb2o_2 _21717_ (.A1_N(_07392_),
    .A2_N(_07396_),
    .B1(_07392_),
    .B2(_07396_),
    .X(_07397_));
 sky130_fd_sc_hd__a2bb2o_2 _21718_ (.A1_N(_07249_),
    .A2_N(_07397_),
    .B1(_07249_),
    .B2(_07397_),
    .X(_07398_));
 sky130_fd_sc_hd__a2bb2o_2 _21719_ (.A1_N(_07391_),
    .A2_N(_07398_),
    .B1(_07391_),
    .B2(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__a2bb2o_2 _21720_ (.A1_N(_07256_),
    .A2_N(_07399_),
    .B1(_07256_),
    .B2(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__a2bb2o_2 _21721_ (.A1_N(_07385_),
    .A2_N(_07400_),
    .B1(_07385_),
    .B2(_07400_),
    .X(_07401_));
 sky130_fd_sc_hd__o22a_2 _21722_ (.A1(_07108_),
    .A2(_07257_),
    .B1(_07245_),
    .B2(_07258_),
    .X(_07402_));
 sky130_fd_sc_hd__a2bb2o_2 _21723_ (.A1_N(_07401_),
    .A2_N(_07402_),
    .B1(_07401_),
    .B2(_07402_),
    .X(_07403_));
 sky130_fd_sc_hd__a2bb2o_2 _21724_ (.A1_N(_07373_),
    .A2_N(_07403_),
    .B1(_07373_),
    .B2(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__o22a_2 _21725_ (.A1(_07119_),
    .A2(_07259_),
    .B1(_07235_),
    .B2(_07260_),
    .X(_07405_));
 sky130_fd_sc_hd__a2bb2o_2 _21726_ (.A1_N(_07404_),
    .A2_N(_07405_),
    .B1(_07404_),
    .B2(_07405_),
    .X(_07406_));
 sky130_fd_sc_hd__a2bb2o_2 _21727_ (.A1_N(_07355_),
    .A2_N(_07406_),
    .B1(_07355_),
    .B2(_07406_),
    .X(_07407_));
 sky130_fd_sc_hd__o22a_2 _21728_ (.A1(_07261_),
    .A2(_07262_),
    .B1(_07218_),
    .B2(_07263_),
    .X(_07408_));
 sky130_fd_sc_hd__a2bb2o_2 _21729_ (.A1_N(_07407_),
    .A2_N(_07408_),
    .B1(_07407_),
    .B2(_07408_),
    .X(_07409_));
 sky130_fd_sc_hd__a2bb2o_2 _21730_ (.A1_N(_07322_),
    .A2_N(_07409_),
    .B1(_07322_),
    .B2(_07409_),
    .X(_07410_));
 sky130_fd_sc_hd__o22a_2 _21731_ (.A1(_07264_),
    .A2(_07265_),
    .B1(_07188_),
    .B2(_07266_),
    .X(_07411_));
 sky130_fd_sc_hd__a2bb2o_2 _21732_ (.A1_N(_07410_),
    .A2_N(_07411_),
    .B1(_07410_),
    .B2(_07411_),
    .X(_07412_));
 sky130_fd_sc_hd__a2bb2o_2 _21733_ (.A1_N(_07281_),
    .A2_N(_07412_),
    .B1(_07281_),
    .B2(_07412_),
    .X(_07413_));
 sky130_fd_sc_hd__o22a_2 _21734_ (.A1(_07267_),
    .A2(_07268_),
    .B1(_07144_),
    .B2(_07269_),
    .X(_07414_));
 sky130_fd_sc_hd__a2bb2o_2 _21735_ (.A1_N(_07413_),
    .A2_N(_07414_),
    .B1(_07413_),
    .B2(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__a2bb2o_2 _21736_ (.A1_N(_07143_),
    .A2_N(_07415_),
    .B1(_07143_),
    .B2(_07415_),
    .X(_07416_));
 sky130_fd_sc_hd__o22a_2 _21737_ (.A1(_07270_),
    .A2(_07271_),
    .B1(_07002_),
    .B2(_07272_),
    .X(_07417_));
 sky130_fd_sc_hd__or2_2 _21738_ (.A(_07416_),
    .B(_07417_),
    .X(_07418_));
 sky130_fd_sc_hd__a21bo_2 _21739_ (.A1(_07416_),
    .A2(_07417_),
    .B1_N(_07418_),
    .X(_07419_));
 sky130_fd_sc_hd__or2_2 _21740_ (.A(_07137_),
    .B(_07276_),
    .X(_07420_));
 sky130_fd_sc_hd__or3_2 _21741_ (.A(_06861_),
    .B(_06998_),
    .C(_07420_),
    .X(_07421_));
 sky130_fd_sc_hd__or2_2 _21742_ (.A(_06863_),
    .B(_07421_),
    .X(_07422_));
 sky130_fd_sc_hd__o221a_2 _21743_ (.A1(_07136_),
    .A2(_07274_),
    .B1(_07138_),
    .B2(_07420_),
    .C1(_07275_),
    .X(_07423_));
 sky130_fd_sc_hd__o21a_2 _21744_ (.A1(_06864_),
    .A2(_07421_),
    .B1(_07423_),
    .X(_07424_));
 sky130_fd_sc_hd__o221a_2 _21745_ (.A1(_06347_),
    .A2(_07422_),
    .B1(_06345_),
    .B2(_07422_),
    .C1(_07424_),
    .X(_07425_));
 sky130_fd_sc_hd__buf_1 _21746_ (.A(_07425_),
    .X(_07426_));
 sky130_fd_sc_hd__a2bb2oi_2 _21747_ (.A1_N(_07419_),
    .A2_N(_07426_),
    .B1(_07419_),
    .B2(_07426_),
    .Y(_02651_));
 sky130_fd_sc_hd__o21ai_2 _21748_ (.A1(_07419_),
    .A2(_07426_),
    .B1(_07418_),
    .Y(_07427_));
 sky130_fd_sc_hd__o22a_2 _21749_ (.A1(_07278_),
    .A2(_07279_),
    .B1(_10600_),
    .B2(_07280_),
    .X(_07428_));
 sky130_fd_sc_hd__o22a_2 _21750_ (.A1(_07283_),
    .A2(_07320_),
    .B1(_07282_),
    .B2(_07321_),
    .X(_07429_));
 sky130_fd_sc_hd__o22a_2 _21751_ (.A1(_07301_),
    .A2(_07302_),
    .B1(_07284_),
    .B2(_07303_),
    .X(_07430_));
 sky130_fd_sc_hd__or2_2 _21752_ (.A(_07429_),
    .B(_07430_),
    .X(_07431_));
 sky130_fd_sc_hd__a21bo_2 _21753_ (.A1(_07429_),
    .A2(_07430_),
    .B1_N(_07431_),
    .X(_07432_));
 sky130_fd_sc_hd__o22a_2 _21754_ (.A1(_07317_),
    .A2(_07318_),
    .B1(_07304_),
    .B2(_07319_),
    .X(_07433_));
 sky130_fd_sc_hd__o22a_2 _21755_ (.A1(_07324_),
    .A2(_07353_),
    .B1(_07323_),
    .B2(_07354_),
    .X(_07434_));
 sky130_fd_sc_hd__a21oi_2 _21756_ (.A1(_07288_),
    .A2(_07290_),
    .B1(_07287_),
    .Y(_07435_));
 sky130_fd_sc_hd__or2_2 _21757_ (.A(_05069_),
    .B(_07159_),
    .X(_07436_));
 sky130_fd_sc_hd__or2_2 _21758_ (.A(_10585_),
    .B(_04693_),
    .X(_07437_));
 sky130_fd_sc_hd__o2bb2a_2 _21759_ (.A1_N(_07436_),
    .A2_N(_07437_),
    .B1(_07436_),
    .B2(_07437_),
    .X(_07438_));
 sky130_vsdinv _21760_ (.A(_07438_),
    .Y(_07439_));
 sky130_fd_sc_hd__or2_2 _21761_ (.A(_05162_),
    .B(_07024_),
    .X(_07440_));
 sky130_fd_sc_hd__a32o_2 _21762_ (.A1(\pcpi_mul.rs2[3] ),
    .A2(_11878_),
    .A3(_07438_),
    .B1(_07439_),
    .B2(_07440_),
    .X(_07441_));
 sky130_fd_sc_hd__o22a_2 _21763_ (.A1(_05171_),
    .A2(_06748_),
    .B1(_05173_),
    .B2(_06890_),
    .X(_07442_));
 sky130_fd_sc_hd__and4_2 _21764_ (.A(_05513_),
    .B(\pcpi_mul.rs1[28] ),
    .C(_05515_),
    .D(\pcpi_mul.rs1[29] ),
    .X(_07443_));
 sky130_fd_sc_hd__or2_2 _21765_ (.A(_07442_),
    .B(_07443_),
    .X(_07444_));
 sky130_vsdinv _21766_ (.A(_07444_),
    .Y(_07445_));
 sky130_fd_sc_hd__a22o_2 _21767_ (.A1(_07297_),
    .A2(_07445_),
    .B1(_07295_),
    .B2(_07444_),
    .X(_07446_));
 sky130_fd_sc_hd__buf_1 _21768_ (.A(_07296_),
    .X(_07447_));
 sky130_fd_sc_hd__a21oi_2 _21769_ (.A1(_07294_),
    .A2(_07447_),
    .B1(_07293_),
    .Y(_07448_));
 sky130_fd_sc_hd__a2bb2o_2 _21770_ (.A1_N(_07446_),
    .A2_N(_07448_),
    .B1(_07446_),
    .B2(_07448_),
    .X(_07449_));
 sky130_fd_sc_hd__a2bb2o_2 _21771_ (.A1_N(_07441_),
    .A2_N(_07449_),
    .B1(_07441_),
    .B2(_07449_),
    .X(_07450_));
 sky130_fd_sc_hd__o22a_2 _21772_ (.A1(_07298_),
    .A2(_07299_),
    .B1(_07291_),
    .B2(_07300_),
    .X(_07451_));
 sky130_fd_sc_hd__a2bb2o_2 _21773_ (.A1_N(_07450_),
    .A2_N(_07451_),
    .B1(_07450_),
    .B2(_07451_),
    .X(_07452_));
 sky130_fd_sc_hd__a2bb2o_2 _21774_ (.A1_N(_07435_),
    .A2_N(_07452_),
    .B1(_07435_),
    .B2(_07452_),
    .X(_07453_));
 sky130_fd_sc_hd__o22a_2 _21775_ (.A1(_07308_),
    .A2(_07313_),
    .B1(_07307_),
    .B2(_07314_),
    .X(_07454_));
 sky130_fd_sc_hd__o22a_2 _21776_ (.A1(_07334_),
    .A2(_07335_),
    .B1(_07329_),
    .B2(_07336_),
    .X(_07455_));
 sky130_fd_sc_hd__a21oi_2 _21777_ (.A1(_07311_),
    .A2(_07312_),
    .B1(_07310_),
    .Y(_07456_));
 sky130_fd_sc_hd__o21ba_2 _21778_ (.A1(_07325_),
    .A2(_07328_),
    .B1_N(_07327_),
    .X(_07457_));
 sky130_fd_sc_hd__o22a_2 _21779_ (.A1(_06132_),
    .A2(_06376_),
    .B1(_06133_),
    .B2(_06742_),
    .X(_07458_));
 sky130_fd_sc_hd__buf_1 _21780_ (.A(\pcpi_mul.rs1[26] ),
    .X(_07459_));
 sky130_fd_sc_hd__and4_2 _21781_ (.A(_06136_),
    .B(_11892_),
    .C(_06137_),
    .D(_07459_),
    .X(_07460_));
 sky130_fd_sc_hd__nor2_2 _21782_ (.A(_07458_),
    .B(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__nor2_2 _21783_ (.A(_04830_),
    .B(_06879_),
    .Y(_07462_));
 sky130_fd_sc_hd__a2bb2o_2 _21784_ (.A1_N(_07461_),
    .A2_N(_07462_),
    .B1(_07461_),
    .B2(_07462_),
    .X(_07463_));
 sky130_fd_sc_hd__a2bb2o_2 _21785_ (.A1_N(_07457_),
    .A2_N(_07463_),
    .B1(_07457_),
    .B2(_07463_),
    .X(_07464_));
 sky130_fd_sc_hd__a2bb2o_2 _21786_ (.A1_N(_07456_),
    .A2_N(_07464_),
    .B1(_07456_),
    .B2(_07464_),
    .X(_07465_));
 sky130_fd_sc_hd__a2bb2o_2 _21787_ (.A1_N(_07455_),
    .A2_N(_07465_),
    .B1(_07455_),
    .B2(_07465_),
    .X(_07466_));
 sky130_fd_sc_hd__a2bb2o_2 _21788_ (.A1_N(_07454_),
    .A2_N(_07466_),
    .B1(_07454_),
    .B2(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__o22a_2 _21789_ (.A1(_07306_),
    .A2(_07315_),
    .B1(_07305_),
    .B2(_07316_),
    .X(_07468_));
 sky130_fd_sc_hd__a2bb2o_2 _21790_ (.A1_N(_07467_),
    .A2_N(_07468_),
    .B1(_07467_),
    .B2(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__a2bb2o_2 _21791_ (.A1_N(_07453_),
    .A2_N(_07469_),
    .B1(_07453_),
    .B2(_07469_),
    .X(_07470_));
 sky130_fd_sc_hd__a2bb2o_2 _21792_ (.A1_N(_07434_),
    .A2_N(_07470_),
    .B1(_07434_),
    .B2(_07470_),
    .X(_07471_));
 sky130_fd_sc_hd__a2bb2o_2 _21793_ (.A1_N(_07433_),
    .A2_N(_07471_),
    .B1(_07433_),
    .B2(_07471_),
    .X(_07472_));
 sky130_fd_sc_hd__o22a_2 _21794_ (.A1(_07350_),
    .A2(_07351_),
    .B1(_07337_),
    .B2(_07352_),
    .X(_07473_));
 sky130_fd_sc_hd__o22a_2 _21795_ (.A1(_07357_),
    .A2(_07371_),
    .B1(_07356_),
    .B2(_07372_),
    .X(_07474_));
 sky130_fd_sc_hd__or2_2 _21796_ (.A(_06049_),
    .B(_06361_),
    .X(_07475_));
 sky130_fd_sc_hd__o22a_2 _21797_ (.A1(_06051_),
    .A2(_05995_),
    .B1(_06052_),
    .B2(_06111_),
    .X(_07476_));
 sky130_fd_sc_hd__and4_2 _21798_ (.A(_06054_),
    .B(_11899_),
    .C(_06055_),
    .D(_07038_),
    .X(_07477_));
 sky130_fd_sc_hd__or2_2 _21799_ (.A(_07476_),
    .B(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__a2bb2o_2 _21800_ (.A1_N(_07475_),
    .A2_N(_07478_),
    .B1(_07475_),
    .B2(_07478_),
    .X(_07479_));
 sky130_fd_sc_hd__or2_2 _21801_ (.A(_06305_),
    .B(_05987_),
    .X(_07480_));
 sky130_fd_sc_hd__buf_1 _21802_ (.A(_05321_),
    .X(_07481_));
 sky130_fd_sc_hd__o22a_2 _21803_ (.A1(_06178_),
    .A2(_05814_),
    .B1(_07481_),
    .B2(_06236_),
    .X(_07482_));
 sky130_fd_sc_hd__buf_1 _21804_ (.A(_11607_),
    .X(_07483_));
 sky130_fd_sc_hd__buf_1 _21805_ (.A(_11610_),
    .X(_07484_));
 sky130_fd_sc_hd__and4_2 _21806_ (.A(_07483_),
    .B(_06517_),
    .C(_07484_),
    .D(_06239_),
    .X(_07485_));
 sky130_fd_sc_hd__or2_2 _21807_ (.A(_07482_),
    .B(_07485_),
    .X(_07486_));
 sky130_fd_sc_hd__a2bb2o_2 _21808_ (.A1_N(_07480_),
    .A2_N(_07486_),
    .B1(_07480_),
    .B2(_07486_),
    .X(_07487_));
 sky130_fd_sc_hd__o21ba_2 _21809_ (.A1(_07330_),
    .A2(_07333_),
    .B1_N(_07332_),
    .X(_07488_));
 sky130_fd_sc_hd__a2bb2o_2 _21810_ (.A1_N(_07487_),
    .A2_N(_07488_),
    .B1(_07487_),
    .B2(_07488_),
    .X(_07489_));
 sky130_fd_sc_hd__a2bb2o_2 _21811_ (.A1_N(_07479_),
    .A2_N(_07489_),
    .B1(_07479_),
    .B2(_07489_),
    .X(_07490_));
 sky130_fd_sc_hd__a21oi_2 _21812_ (.A1(_07345_),
    .A2(_07347_),
    .B1(_07344_),
    .Y(_07491_));
 sky130_fd_sc_hd__o21ba_2 _21813_ (.A1(_07358_),
    .A2(_07362_),
    .B1_N(_07361_),
    .X(_07492_));
 sky130_fd_sc_hd__or2_2 _21814_ (.A(_05309_),
    .B(_06255_),
    .X(_07493_));
 sky130_fd_sc_hd__o22a_2 _21815_ (.A1(_07340_),
    .A2(_05501_),
    .B1(_06549_),
    .B2(_06257_),
    .X(_07494_));
 sky130_fd_sc_hd__and4_2 _21816_ (.A(_07342_),
    .B(_06138_),
    .C(_07343_),
    .D(_06392_),
    .X(_07495_));
 sky130_fd_sc_hd__or2_2 _21817_ (.A(_07494_),
    .B(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__a2bb2o_2 _21818_ (.A1_N(_07493_),
    .A2_N(_07496_),
    .B1(_07493_),
    .B2(_07496_),
    .X(_07497_));
 sky130_fd_sc_hd__a2bb2o_2 _21819_ (.A1_N(_07492_),
    .A2_N(_07497_),
    .B1(_07492_),
    .B2(_07497_),
    .X(_07498_));
 sky130_fd_sc_hd__a2bb2o_2 _21820_ (.A1_N(_07491_),
    .A2_N(_07498_),
    .B1(_07491_),
    .B2(_07498_),
    .X(_07499_));
 sky130_fd_sc_hd__o22a_2 _21821_ (.A1(_07339_),
    .A2(_07348_),
    .B1(_07338_),
    .B2(_07349_),
    .X(_07500_));
 sky130_fd_sc_hd__a2bb2o_2 _21822_ (.A1_N(_07499_),
    .A2_N(_07500_),
    .B1(_07499_),
    .B2(_07500_),
    .X(_07501_));
 sky130_fd_sc_hd__a2bb2o_2 _21823_ (.A1_N(_07490_),
    .A2_N(_07501_),
    .B1(_07490_),
    .B2(_07501_),
    .X(_07502_));
 sky130_fd_sc_hd__a2bb2o_2 _21824_ (.A1_N(_07474_),
    .A2_N(_07502_),
    .B1(_07474_),
    .B2(_07502_),
    .X(_07503_));
 sky130_fd_sc_hd__a2bb2o_2 _21825_ (.A1_N(_07473_),
    .A2_N(_07503_),
    .B1(_07473_),
    .B2(_07503_),
    .X(_07504_));
 sky130_fd_sc_hd__o22a_2 _21826_ (.A1(_07368_),
    .A2(_07369_),
    .B1(_07363_),
    .B2(_07370_),
    .X(_07505_));
 sky130_fd_sc_hd__o22a_2 _21827_ (.A1(_07375_),
    .A2(_07383_),
    .B1(_07374_),
    .B2(_07384_),
    .X(_07506_));
 sky130_fd_sc_hd__or2_2 _21828_ (.A(_06700_),
    .B(_05720_),
    .X(_07507_));
 sky130_fd_sc_hd__o22a_2 _21829_ (.A1(_07359_),
    .A2(_05609_),
    .B1(_05662_),
    .B2(_05334_),
    .X(_07508_));
 sky130_fd_sc_hd__buf_1 _21830_ (.A(\pcpi_mul.rs1[14] ),
    .X(_07509_));
 sky130_fd_sc_hd__and4_2 _21831_ (.A(_06703_),
    .B(_05848_),
    .C(_06570_),
    .D(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__or2_2 _21832_ (.A(_07508_),
    .B(_07510_),
    .X(_07511_));
 sky130_fd_sc_hd__a2bb2o_2 _21833_ (.A1_N(_07507_),
    .A2_N(_07511_),
    .B1(_07507_),
    .B2(_07511_),
    .X(_07512_));
 sky130_fd_sc_hd__or2_2 _21834_ (.A(_05926_),
    .B(_05158_),
    .X(_07513_));
 sky130_fd_sc_hd__o22a_2 _21835_ (.A1(_06818_),
    .A2(_06180_),
    .B1(_06030_),
    .B2(_05530_),
    .X(_07514_));
 sky130_fd_sc_hd__buf_1 _21836_ (.A(_11584_),
    .X(_07515_));
 sky130_fd_sc_hd__buf_1 _21837_ (.A(_11588_),
    .X(_07516_));
 sky130_fd_sc_hd__and4_2 _21838_ (.A(_07515_),
    .B(_11929_),
    .C(_07516_),
    .D(_05743_),
    .X(_07517_));
 sky130_fd_sc_hd__or2_2 _21839_ (.A(_07514_),
    .B(_07517_),
    .X(_07518_));
 sky130_fd_sc_hd__a2bb2o_2 _21840_ (.A1_N(_07513_),
    .A2_N(_07518_),
    .B1(_07513_),
    .B2(_07518_),
    .X(_07519_));
 sky130_fd_sc_hd__o21ba_2 _21841_ (.A1(_07364_),
    .A2(_07367_),
    .B1_N(_07366_),
    .X(_07520_));
 sky130_fd_sc_hd__a2bb2o_2 _21842_ (.A1_N(_07519_),
    .A2_N(_07520_),
    .B1(_07519_),
    .B2(_07520_),
    .X(_07521_));
 sky130_fd_sc_hd__a2bb2o_2 _21843_ (.A1_N(_07512_),
    .A2_N(_07521_),
    .B1(_07512_),
    .B2(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__a2bb2o_2 _21844_ (.A1_N(_07506_),
    .A2_N(_07522_),
    .B1(_07506_),
    .B2(_07522_),
    .X(_07523_));
 sky130_fd_sc_hd__a2bb2o_2 _21845_ (.A1_N(_07505_),
    .A2_N(_07523_),
    .B1(_07505_),
    .B2(_07523_),
    .X(_07524_));
 sky130_fd_sc_hd__o21ba_2 _21846_ (.A1(_07377_),
    .A2(_07382_),
    .B1_N(_07381_),
    .X(_07525_));
 sky130_fd_sc_hd__o21ba_2 _21847_ (.A1(_07386_),
    .A2(_07390_),
    .B1_N(_07389_),
    .X(_07526_));
 sky130_fd_sc_hd__or2_2 _21848_ (.A(_07376_),
    .B(_05077_),
    .X(_07527_));
 sky130_fd_sc_hd__o22a_2 _21849_ (.A1(_07378_),
    .A2(_05396_),
    .B1(_07379_),
    .B2(_06568_),
    .X(_07528_));
 sky130_fd_sc_hd__and4_2 _21850_ (.A(_07240_),
    .B(_11937_),
    .C(_11580_),
    .D(_11934_),
    .X(_07529_));
 sky130_fd_sc_hd__or2_2 _21851_ (.A(_07528_),
    .B(_07529_),
    .X(_07530_));
 sky130_fd_sc_hd__a2bb2o_2 _21852_ (.A1_N(_07527_),
    .A2_N(_07530_),
    .B1(_07527_),
    .B2(_07530_),
    .X(_07531_));
 sky130_fd_sc_hd__a2bb2o_2 _21853_ (.A1_N(_07526_),
    .A2_N(_07531_),
    .B1(_07526_),
    .B2(_07531_),
    .X(_07532_));
 sky130_fd_sc_hd__a2bb2o_2 _21854_ (.A1_N(_07525_),
    .A2_N(_07532_),
    .B1(_07525_),
    .B2(_07532_),
    .X(_07533_));
 sky130_fd_sc_hd__or2_2 _21855_ (.A(_06685_),
    .B(_06277_),
    .X(_07534_));
 sky130_fd_sc_hd__buf_1 _21856_ (.A(_07387_),
    .X(_07535_));
 sky130_fd_sc_hd__buf_1 _21857_ (.A(_06829_),
    .X(_07536_));
 sky130_fd_sc_hd__o22a_2 _21858_ (.A1(_07535_),
    .A2(_05403_),
    .B1(_07536_),
    .B2(_06151_),
    .X(_07537_));
 sky130_fd_sc_hd__buf_1 _21859_ (.A(_11566_),
    .X(_07538_));
 sky130_fd_sc_hd__buf_1 _21860_ (.A(_11570_),
    .X(_07539_));
 sky130_fd_sc_hd__and4_2 _21861_ (.A(_07538_),
    .B(_11946_),
    .C(_07539_),
    .D(_11943_),
    .X(_07540_));
 sky130_fd_sc_hd__or2_2 _21862_ (.A(_07537_),
    .B(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__a2bb2o_2 _21863_ (.A1_N(_07534_),
    .A2_N(_07541_),
    .B1(_07534_),
    .B2(_07541_),
    .X(_07542_));
 sky130_fd_sc_hd__or2_2 _21864_ (.A(_07100_),
    .B(_04723_),
    .X(_07543_));
 sky130_fd_sc_hd__and4_2 _21865_ (.A(_07393_),
    .B(_04709_),
    .C(_11559_),
    .D(_11952_),
    .X(_07544_));
 sky130_fd_sc_hd__buf_1 _21866_ (.A(_07246_),
    .X(_07545_));
 sky130_fd_sc_hd__o22a_2 _21867_ (.A1(_10596_),
    .A2(_11955_),
    .B1(_07545_),
    .B2(_05061_),
    .X(_07546_));
 sky130_fd_sc_hd__or2_2 _21868_ (.A(_07544_),
    .B(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__a2bb2o_2 _21869_ (.A1_N(_07543_),
    .A2_N(_07547_),
    .B1(_07543_),
    .B2(_07547_),
    .X(_07548_));
 sky130_fd_sc_hd__o21ba_2 _21870_ (.A1(_07392_),
    .A2(_07396_),
    .B1_N(_07394_),
    .X(_07549_));
 sky130_fd_sc_hd__a2bb2o_2 _21871_ (.A1_N(_07548_),
    .A2_N(_07549_),
    .B1(_07548_),
    .B2(_07549_),
    .X(_07550_));
 sky130_fd_sc_hd__a2bb2o_2 _21872_ (.A1_N(_07542_),
    .A2_N(_07550_),
    .B1(_07542_),
    .B2(_07550_),
    .X(_07551_));
 sky130_fd_sc_hd__o22a_2 _21873_ (.A1(_07249_),
    .A2(_07397_),
    .B1(_07391_),
    .B2(_07398_),
    .X(_07552_));
 sky130_fd_sc_hd__a2bb2o_2 _21874_ (.A1_N(_07551_),
    .A2_N(_07552_),
    .B1(_07551_),
    .B2(_07552_),
    .X(_07553_));
 sky130_fd_sc_hd__a2bb2o_2 _21875_ (.A1_N(_07533_),
    .A2_N(_07553_),
    .B1(_07533_),
    .B2(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__o22a_2 _21876_ (.A1(_07256_),
    .A2(_07399_),
    .B1(_07385_),
    .B2(_07400_),
    .X(_07555_));
 sky130_fd_sc_hd__a2bb2o_2 _21877_ (.A1_N(_07554_),
    .A2_N(_07555_),
    .B1(_07554_),
    .B2(_07555_),
    .X(_07556_));
 sky130_fd_sc_hd__a2bb2o_2 _21878_ (.A1_N(_07524_),
    .A2_N(_07556_),
    .B1(_07524_),
    .B2(_07556_),
    .X(_07557_));
 sky130_fd_sc_hd__o22a_2 _21879_ (.A1(_07401_),
    .A2(_07402_),
    .B1(_07373_),
    .B2(_07403_),
    .X(_07558_));
 sky130_fd_sc_hd__a2bb2o_2 _21880_ (.A1_N(_07557_),
    .A2_N(_07558_),
    .B1(_07557_),
    .B2(_07558_),
    .X(_07559_));
 sky130_fd_sc_hd__a2bb2o_2 _21881_ (.A1_N(_07504_),
    .A2_N(_07559_),
    .B1(_07504_),
    .B2(_07559_),
    .X(_07560_));
 sky130_fd_sc_hd__o22a_2 _21882_ (.A1(_07404_),
    .A2(_07405_),
    .B1(_07355_),
    .B2(_07406_),
    .X(_07561_));
 sky130_fd_sc_hd__a2bb2o_2 _21883_ (.A1_N(_07560_),
    .A2_N(_07561_),
    .B1(_07560_),
    .B2(_07561_),
    .X(_07562_));
 sky130_fd_sc_hd__a2bb2o_2 _21884_ (.A1_N(_07472_),
    .A2_N(_07562_),
    .B1(_07472_),
    .B2(_07562_),
    .X(_07563_));
 sky130_fd_sc_hd__o22a_2 _21885_ (.A1(_07407_),
    .A2(_07408_),
    .B1(_07322_),
    .B2(_07409_),
    .X(_07564_));
 sky130_fd_sc_hd__a2bb2o_2 _21886_ (.A1_N(_07563_),
    .A2_N(_07564_),
    .B1(_07563_),
    .B2(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__a2bb2o_2 _21887_ (.A1_N(_07432_),
    .A2_N(_07565_),
    .B1(_07432_),
    .B2(_07565_),
    .X(_07566_));
 sky130_fd_sc_hd__o22a_2 _21888_ (.A1(_07410_),
    .A2(_07411_),
    .B1(_07281_),
    .B2(_07412_),
    .X(_07567_));
 sky130_fd_sc_hd__a2bb2o_2 _21889_ (.A1_N(_07566_),
    .A2_N(_07567_),
    .B1(_07566_),
    .B2(_07567_),
    .X(_07568_));
 sky130_fd_sc_hd__a2bb2o_2 _21890_ (.A1_N(_07428_),
    .A2_N(_07568_),
    .B1(_07428_),
    .B2(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__o22a_2 _21891_ (.A1(_07413_),
    .A2(_07414_),
    .B1(_07143_),
    .B2(_07415_),
    .X(_07570_));
 sky130_fd_sc_hd__or2_2 _21892_ (.A(_07569_),
    .B(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__a21bo_2 _21893_ (.A1(_07569_),
    .A2(_07570_),
    .B1_N(_07571_),
    .X(_07572_));
 sky130_fd_sc_hd__a2bb2o_2 _21894_ (.A1_N(_07427_),
    .A2_N(_07572_),
    .B1(_07427_),
    .B2(_07572_),
    .X(_02652_));
 sky130_fd_sc_hd__o22a_2 _21895_ (.A1(_07434_),
    .A2(_07470_),
    .B1(_07433_),
    .B2(_07471_),
    .X(_07573_));
 sky130_fd_sc_hd__o22a_2 _21896_ (.A1(_07450_),
    .A2(_07451_),
    .B1(_07435_),
    .B2(_07452_),
    .X(_07574_));
 sky130_fd_sc_hd__or2_2 _21897_ (.A(_07573_),
    .B(_07574_),
    .X(_07575_));
 sky130_fd_sc_hd__a21bo_2 _21898_ (.A1(_07573_),
    .A2(_07574_),
    .B1_N(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__o22a_2 _21899_ (.A1(_07467_),
    .A2(_07468_),
    .B1(_07453_),
    .B2(_07469_),
    .X(_07577_));
 sky130_fd_sc_hd__o22a_2 _21900_ (.A1(_07474_),
    .A2(_07502_),
    .B1(_07473_),
    .B2(_07503_),
    .X(_07578_));
 sky130_fd_sc_hd__o22a_2 _21901_ (.A1(_07436_),
    .A2(_07437_),
    .B1(_07439_),
    .B2(_07440_),
    .X(_07579_));
 sky130_fd_sc_hd__or2_2 _21902_ (.A(_10585_),
    .B(_04706_),
    .X(_07580_));
 sky130_fd_sc_hd__nor2_2 _21903_ (.A(_07437_),
    .B(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__a21oi_2 _21904_ (.A1(_07437_),
    .A2(_07580_),
    .B1(_07581_),
    .Y(_07582_));
 sky130_fd_sc_hd__buf_1 _21905_ (.A(_07160_),
    .X(_07583_));
 sky130_fd_sc_hd__nor2_2 _21906_ (.A(_06107_),
    .B(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__a2bb2o_2 _21907_ (.A1_N(_07582_),
    .A2_N(_07584_),
    .B1(_07582_),
    .B2(_07584_),
    .X(_07585_));
 sky130_fd_sc_hd__o22a_2 _21908_ (.A1(_05826_),
    .A2(_06890_),
    .B1(_05827_),
    .B2(_07022_),
    .X(_07586_));
 sky130_fd_sc_hd__buf_1 _21909_ (.A(\pcpi_mul.rs1[29] ),
    .X(_07587_));
 sky130_fd_sc_hd__and4_2 _21910_ (.A(_05513_),
    .B(_07587_),
    .C(_05515_),
    .D(_11876_),
    .X(_07588_));
 sky130_fd_sc_hd__or2_2 _21911_ (.A(_07586_),
    .B(_07588_),
    .X(_07589_));
 sky130_vsdinv _21912_ (.A(_07589_),
    .Y(_07590_));
 sky130_fd_sc_hd__a22o_2 _21913_ (.A1(_07297_),
    .A2(_07590_),
    .B1(_07295_),
    .B2(_07589_),
    .X(_07591_));
 sky130_fd_sc_hd__a21oi_2 _21914_ (.A1(_07447_),
    .A2(_07445_),
    .B1(_07443_),
    .Y(_07592_));
 sky130_fd_sc_hd__a2bb2o_2 _21915_ (.A1_N(_07591_),
    .A2_N(_07592_),
    .B1(_07591_),
    .B2(_07592_),
    .X(_07593_));
 sky130_fd_sc_hd__a2bb2o_2 _21916_ (.A1_N(_07585_),
    .A2_N(_07593_),
    .B1(_07585_),
    .B2(_07593_),
    .X(_07594_));
 sky130_fd_sc_hd__o22a_2 _21917_ (.A1(_07446_),
    .A2(_07448_),
    .B1(_07441_),
    .B2(_07449_),
    .X(_07595_));
 sky130_fd_sc_hd__a2bb2o_2 _21918_ (.A1_N(_07594_),
    .A2_N(_07595_),
    .B1(_07594_),
    .B2(_07595_),
    .X(_07596_));
 sky130_fd_sc_hd__a2bb2o_2 _21919_ (.A1_N(_07579_),
    .A2_N(_07596_),
    .B1(_07579_),
    .B2(_07596_),
    .X(_07597_));
 sky130_fd_sc_hd__o22a_2 _21920_ (.A1(_07457_),
    .A2(_07463_),
    .B1(_07456_),
    .B2(_07464_),
    .X(_07598_));
 sky130_fd_sc_hd__o22a_2 _21921_ (.A1(_07487_),
    .A2(_07488_),
    .B1(_07479_),
    .B2(_07489_),
    .X(_07599_));
 sky130_fd_sc_hd__a21oi_2 _21922_ (.A1(_07461_),
    .A2(_07462_),
    .B1(_07460_),
    .Y(_07600_));
 sky130_fd_sc_hd__o21ba_2 _21923_ (.A1(_07475_),
    .A2(_07478_),
    .B1_N(_07477_),
    .X(_07601_));
 sky130_fd_sc_hd__buf_1 _21924_ (.A(_05193_),
    .X(_07602_));
 sky130_fd_sc_hd__o22a_2 _21925_ (.A1(_07602_),
    .A2(_06742_),
    .B1(_04828_),
    .B2(_06878_),
    .X(_07603_));
 sky130_fd_sc_hd__and4_2 _21926_ (.A(_11620_),
    .B(_07459_),
    .C(_11624_),
    .D(_11884_),
    .X(_07604_));
 sky130_fd_sc_hd__nor2_2 _21927_ (.A(_07603_),
    .B(_07604_),
    .Y(_07605_));
 sky130_fd_sc_hd__nor2_2 _21928_ (.A(_04795_),
    .B(_06750_),
    .Y(_07606_));
 sky130_fd_sc_hd__a2bb2o_2 _21929_ (.A1_N(_07605_),
    .A2_N(_07606_),
    .B1(_07605_),
    .B2(_07606_),
    .X(_07607_));
 sky130_fd_sc_hd__a2bb2o_2 _21930_ (.A1_N(_07601_),
    .A2_N(_07607_),
    .B1(_07601_),
    .B2(_07607_),
    .X(_07608_));
 sky130_fd_sc_hd__a2bb2o_2 _21931_ (.A1_N(_07600_),
    .A2_N(_07608_),
    .B1(_07600_),
    .B2(_07608_),
    .X(_07609_));
 sky130_fd_sc_hd__a2bb2o_2 _21932_ (.A1_N(_07599_),
    .A2_N(_07609_),
    .B1(_07599_),
    .B2(_07609_),
    .X(_07610_));
 sky130_fd_sc_hd__a2bb2o_2 _21933_ (.A1_N(_07598_),
    .A2_N(_07610_),
    .B1(_07598_),
    .B2(_07610_),
    .X(_07611_));
 sky130_fd_sc_hd__o22a_2 _21934_ (.A1(_07455_),
    .A2(_07465_),
    .B1(_07454_),
    .B2(_07466_),
    .X(_07612_));
 sky130_fd_sc_hd__a2bb2o_2 _21935_ (.A1_N(_07611_),
    .A2_N(_07612_),
    .B1(_07611_),
    .B2(_07612_),
    .X(_07613_));
 sky130_fd_sc_hd__a2bb2o_2 _21936_ (.A1_N(_07597_),
    .A2_N(_07613_),
    .B1(_07597_),
    .B2(_07613_),
    .X(_07614_));
 sky130_fd_sc_hd__a2bb2o_2 _21937_ (.A1_N(_07578_),
    .A2_N(_07614_),
    .B1(_07578_),
    .B2(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__a2bb2o_2 _21938_ (.A1_N(_07577_),
    .A2_N(_07615_),
    .B1(_07577_),
    .B2(_07615_),
    .X(_07616_));
 sky130_fd_sc_hd__o22a_2 _21939_ (.A1(_07499_),
    .A2(_07500_),
    .B1(_07490_),
    .B2(_07501_),
    .X(_07617_));
 sky130_fd_sc_hd__o22a_2 _21940_ (.A1(_07506_),
    .A2(_07522_),
    .B1(_07505_),
    .B2(_07523_),
    .X(_07618_));
 sky130_fd_sc_hd__or2_2 _21941_ (.A(_06049_),
    .B(_06377_),
    .X(_07619_));
 sky130_fd_sc_hd__o22a_2 _21942_ (.A1(_06051_),
    .A2(_06111_),
    .B1(_06052_),
    .B2(_07173_),
    .X(_07620_));
 sky130_fd_sc_hd__and4_2 _21943_ (.A(_06054_),
    .B(_07038_),
    .C(_06055_),
    .D(_07175_),
    .X(_07621_));
 sky130_fd_sc_hd__or2_2 _21944_ (.A(_07620_),
    .B(_07621_),
    .X(_07622_));
 sky130_fd_sc_hd__a2bb2o_2 _21945_ (.A1_N(_07619_),
    .A2_N(_07622_),
    .B1(_07619_),
    .B2(_07622_),
    .X(_07623_));
 sky130_fd_sc_hd__buf_1 _21946_ (.A(_05056_),
    .X(_07624_));
 sky130_fd_sc_hd__or2_2 _21947_ (.A(_07624_),
    .B(_05996_),
    .X(_07625_));
 sky130_fd_sc_hd__buf_1 _21948_ (.A(_05405_),
    .X(_07626_));
 sky130_fd_sc_hd__o22a_2 _21949_ (.A1(_07626_),
    .A2(_05823_),
    .B1(_07481_),
    .B2(_05986_),
    .X(_07627_));
 sky130_fd_sc_hd__and4_2 _21950_ (.A(_07483_),
    .B(_11905_),
    .C(_07484_),
    .D(_06371_),
    .X(_07628_));
 sky130_fd_sc_hd__or2_2 _21951_ (.A(_07627_),
    .B(_07628_),
    .X(_07629_));
 sky130_fd_sc_hd__a2bb2o_2 _21952_ (.A1_N(_07625_),
    .A2_N(_07629_),
    .B1(_07625_),
    .B2(_07629_),
    .X(_07630_));
 sky130_fd_sc_hd__o21ba_2 _21953_ (.A1(_07480_),
    .A2(_07486_),
    .B1_N(_07485_),
    .X(_07631_));
 sky130_fd_sc_hd__a2bb2o_2 _21954_ (.A1_N(_07630_),
    .A2_N(_07631_),
    .B1(_07630_),
    .B2(_07631_),
    .X(_07632_));
 sky130_fd_sc_hd__a2bb2o_2 _21955_ (.A1_N(_07623_),
    .A2_N(_07632_),
    .B1(_07623_),
    .B2(_07632_),
    .X(_07633_));
 sky130_fd_sc_hd__o21ba_2 _21956_ (.A1(_07493_),
    .A2(_07496_),
    .B1_N(_07495_),
    .X(_07634_));
 sky130_fd_sc_hd__o21ba_2 _21957_ (.A1(_07507_),
    .A2(_07511_),
    .B1_N(_07510_),
    .X(_07635_));
 sky130_fd_sc_hd__or2_2 _21958_ (.A(_07346_),
    .B(_05716_),
    .X(_07636_));
 sky130_fd_sc_hd__o22a_2 _21959_ (.A1(_07340_),
    .A2(_06257_),
    .B1(_06549_),
    .B2(_06254_),
    .X(_07637_));
 sky130_fd_sc_hd__and4_2 _21960_ (.A(_07342_),
    .B(_06392_),
    .C(_07343_),
    .D(_06393_),
    .X(_07638_));
 sky130_fd_sc_hd__or2_2 _21961_ (.A(_07637_),
    .B(_07638_),
    .X(_07639_));
 sky130_fd_sc_hd__a2bb2o_2 _21962_ (.A1_N(_07636_),
    .A2_N(_07639_),
    .B1(_07636_),
    .B2(_07639_),
    .X(_07640_));
 sky130_fd_sc_hd__a2bb2o_2 _21963_ (.A1_N(_07635_),
    .A2_N(_07640_),
    .B1(_07635_),
    .B2(_07640_),
    .X(_07641_));
 sky130_fd_sc_hd__a2bb2o_2 _21964_ (.A1_N(_07634_),
    .A2_N(_07641_),
    .B1(_07634_),
    .B2(_07641_),
    .X(_07642_));
 sky130_fd_sc_hd__o22a_2 _21965_ (.A1(_07492_),
    .A2(_07497_),
    .B1(_07491_),
    .B2(_07498_),
    .X(_07643_));
 sky130_fd_sc_hd__a2bb2o_2 _21966_ (.A1_N(_07642_),
    .A2_N(_07643_),
    .B1(_07642_),
    .B2(_07643_),
    .X(_07644_));
 sky130_fd_sc_hd__a2bb2o_2 _21967_ (.A1_N(_07633_),
    .A2_N(_07644_),
    .B1(_07633_),
    .B2(_07644_),
    .X(_07645_));
 sky130_fd_sc_hd__a2bb2o_2 _21968_ (.A1_N(_07618_),
    .A2_N(_07645_),
    .B1(_07618_),
    .B2(_07645_),
    .X(_07646_));
 sky130_fd_sc_hd__a2bb2o_2 _21969_ (.A1_N(_07617_),
    .A2_N(_07646_),
    .B1(_07617_),
    .B2(_07646_),
    .X(_07647_));
 sky130_fd_sc_hd__o22a_2 _21970_ (.A1(_07519_),
    .A2(_07520_),
    .B1(_07512_),
    .B2(_07521_),
    .X(_07648_));
 sky130_fd_sc_hd__o22a_2 _21971_ (.A1(_07526_),
    .A2(_07531_),
    .B1(_07525_),
    .B2(_07532_),
    .X(_07649_));
 sky130_fd_sc_hd__or2_2 _21972_ (.A(_05562_),
    .B(_05502_),
    .X(_07650_));
 sky130_fd_sc_hd__buf_1 _21973_ (.A(_06039_),
    .X(_07651_));
 sky130_fd_sc_hd__o22a_2 _21974_ (.A1(_07651_),
    .A2(_05334_),
    .B1(_05659_),
    .B2(_05420_),
    .X(_07652_));
 sky130_fd_sc_hd__and4_2 _21975_ (.A(_11593_),
    .B(_07509_),
    .C(_11598_),
    .D(_05830_),
    .X(_07653_));
 sky130_fd_sc_hd__or2_2 _21976_ (.A(_07652_),
    .B(_07653_),
    .X(_07654_));
 sky130_fd_sc_hd__a2bb2o_2 _21977_ (.A1_N(_07650_),
    .A2_N(_07654_),
    .B1(_07650_),
    .B2(_07654_),
    .X(_07655_));
 sky130_fd_sc_hd__buf_1 _21978_ (.A(_06035_),
    .X(_07656_));
 sky130_fd_sc_hd__or2_2 _21979_ (.A(_07656_),
    .B(_05247_),
    .X(_07657_));
 sky130_fd_sc_hd__buf_1 _21980_ (.A(_06579_),
    .X(_07658_));
 sky130_fd_sc_hd__o22a_2 _21981_ (.A1(_07658_),
    .A2(_05530_),
    .B1(_06034_),
    .B2(_05740_),
    .X(_07659_));
 sky130_fd_sc_hd__and4_2 _21982_ (.A(_07515_),
    .B(_11927_),
    .C(_07516_),
    .D(_11925_),
    .X(_07660_));
 sky130_fd_sc_hd__or2_2 _21983_ (.A(_07659_),
    .B(_07660_),
    .X(_07661_));
 sky130_fd_sc_hd__a2bb2o_2 _21984_ (.A1_N(_07657_),
    .A2_N(_07661_),
    .B1(_07657_),
    .B2(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__o21ba_2 _21985_ (.A1(_07513_),
    .A2(_07518_),
    .B1_N(_07517_),
    .X(_07663_));
 sky130_fd_sc_hd__a2bb2o_2 _21986_ (.A1_N(_07662_),
    .A2_N(_07663_),
    .B1(_07662_),
    .B2(_07663_),
    .X(_07664_));
 sky130_fd_sc_hd__a2bb2o_2 _21987_ (.A1_N(_07655_),
    .A2_N(_07664_),
    .B1(_07655_),
    .B2(_07664_),
    .X(_07665_));
 sky130_fd_sc_hd__a2bb2o_2 _21988_ (.A1_N(_07649_),
    .A2_N(_07665_),
    .B1(_07649_),
    .B2(_07665_),
    .X(_07666_));
 sky130_fd_sc_hd__a2bb2o_2 _21989_ (.A1_N(_07648_),
    .A2_N(_07666_),
    .B1(_07648_),
    .B2(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__o21ba_2 _21990_ (.A1(_07527_),
    .A2(_07530_),
    .B1_N(_07529_),
    .X(_07668_));
 sky130_fd_sc_hd__o21ba_2 _21991_ (.A1(_07534_),
    .A2(_07541_),
    .B1_N(_07540_),
    .X(_07669_));
 sky130_fd_sc_hd__or2_2 _21992_ (.A(_07376_),
    .B(_05164_),
    .X(_07670_));
 sky130_fd_sc_hd__o22a_2 _21993_ (.A1(_07378_),
    .A2(_05017_),
    .B1(_07379_),
    .B2(_05943_),
    .X(_07671_));
 sky130_fd_sc_hd__buf_1 _21994_ (.A(_11579_),
    .X(_07672_));
 sky130_fd_sc_hd__and4_2 _21995_ (.A(_07240_),
    .B(_11934_),
    .C(_07672_),
    .D(_11931_),
    .X(_07673_));
 sky130_fd_sc_hd__or2_2 _21996_ (.A(_07671_),
    .B(_07673_),
    .X(_07674_));
 sky130_fd_sc_hd__a2bb2o_2 _21997_ (.A1_N(_07670_),
    .A2_N(_07674_),
    .B1(_07670_),
    .B2(_07674_),
    .X(_07675_));
 sky130_fd_sc_hd__a2bb2o_2 _21998_ (.A1_N(_07669_),
    .A2_N(_07675_),
    .B1(_07669_),
    .B2(_07675_),
    .X(_07676_));
 sky130_fd_sc_hd__a2bb2o_2 _21999_ (.A1_N(_07668_),
    .A2_N(_07676_),
    .B1(_07668_),
    .B2(_07676_),
    .X(_07677_));
 sky130_fd_sc_hd__or2_2 _22000_ (.A(_06686_),
    .B(_05191_),
    .X(_07678_));
 sky130_fd_sc_hd__o22a_2 _22001_ (.A1(_07535_),
    .A2(_06151_),
    .B1(_07536_),
    .B2(_06277_),
    .X(_07679_));
 sky130_fd_sc_hd__buf_1 _22002_ (.A(_11566_),
    .X(_07680_));
 sky130_fd_sc_hd__buf_1 _22003_ (.A(_11570_),
    .X(_07681_));
 sky130_fd_sc_hd__and4_2 _22004_ (.A(_07680_),
    .B(_11943_),
    .C(_07681_),
    .D(_11940_),
    .X(_07682_));
 sky130_fd_sc_hd__or2_2 _22005_ (.A(_07679_),
    .B(_07682_),
    .X(_07683_));
 sky130_fd_sc_hd__a2bb2o_2 _22006_ (.A1_N(_07678_),
    .A2_N(_07683_),
    .B1(_07678_),
    .B2(_07683_),
    .X(_07684_));
 sky130_fd_sc_hd__or2_2 _22007_ (.A(_07100_),
    .B(_05403_),
    .X(_07685_));
 sky130_fd_sc_hd__buf_1 _22008_ (.A(_07393_),
    .X(_07686_));
 sky130_fd_sc_hd__and4_2 _22009_ (.A(_07686_),
    .B(_04779_),
    .C(_11559_),
    .D(_11949_),
    .X(_07687_));
 sky130_fd_sc_hd__o22a_2 _22010_ (.A1(_10596_),
    .A2(_11952_),
    .B1(_07545_),
    .B2(_05406_),
    .X(_07688_));
 sky130_fd_sc_hd__or2_2 _22011_ (.A(_07687_),
    .B(_07688_),
    .X(_07689_));
 sky130_fd_sc_hd__a2bb2o_2 _22012_ (.A1_N(_07685_),
    .A2_N(_07689_),
    .B1(_07685_),
    .B2(_07689_),
    .X(_07690_));
 sky130_fd_sc_hd__o21ba_2 _22013_ (.A1(_07543_),
    .A2(_07547_),
    .B1_N(_07544_),
    .X(_07691_));
 sky130_fd_sc_hd__a2bb2o_2 _22014_ (.A1_N(_07690_),
    .A2_N(_07691_),
    .B1(_07690_),
    .B2(_07691_),
    .X(_07692_));
 sky130_fd_sc_hd__a2bb2o_2 _22015_ (.A1_N(_07684_),
    .A2_N(_07692_),
    .B1(_07684_),
    .B2(_07692_),
    .X(_07693_));
 sky130_fd_sc_hd__o22a_2 _22016_ (.A1(_07548_),
    .A2(_07549_),
    .B1(_07542_),
    .B2(_07550_),
    .X(_07694_));
 sky130_fd_sc_hd__a2bb2o_2 _22017_ (.A1_N(_07693_),
    .A2_N(_07694_),
    .B1(_07693_),
    .B2(_07694_),
    .X(_07695_));
 sky130_fd_sc_hd__a2bb2o_2 _22018_ (.A1_N(_07677_),
    .A2_N(_07695_),
    .B1(_07677_),
    .B2(_07695_),
    .X(_07696_));
 sky130_fd_sc_hd__o22a_2 _22019_ (.A1(_07551_),
    .A2(_07552_),
    .B1(_07533_),
    .B2(_07553_),
    .X(_07697_));
 sky130_fd_sc_hd__a2bb2o_2 _22020_ (.A1_N(_07696_),
    .A2_N(_07697_),
    .B1(_07696_),
    .B2(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__a2bb2o_2 _22021_ (.A1_N(_07667_),
    .A2_N(_07698_),
    .B1(_07667_),
    .B2(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__o22a_2 _22022_ (.A1(_07554_),
    .A2(_07555_),
    .B1(_07524_),
    .B2(_07556_),
    .X(_07700_));
 sky130_fd_sc_hd__a2bb2o_2 _22023_ (.A1_N(_07699_),
    .A2_N(_07700_),
    .B1(_07699_),
    .B2(_07700_),
    .X(_07701_));
 sky130_fd_sc_hd__a2bb2o_2 _22024_ (.A1_N(_07647_),
    .A2_N(_07701_),
    .B1(_07647_),
    .B2(_07701_),
    .X(_07702_));
 sky130_fd_sc_hd__o22a_2 _22025_ (.A1(_07557_),
    .A2(_07558_),
    .B1(_07504_),
    .B2(_07559_),
    .X(_07703_));
 sky130_fd_sc_hd__a2bb2o_2 _22026_ (.A1_N(_07702_),
    .A2_N(_07703_),
    .B1(_07702_),
    .B2(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__a2bb2o_2 _22027_ (.A1_N(_07616_),
    .A2_N(_07704_),
    .B1(_07616_),
    .B2(_07704_),
    .X(_07705_));
 sky130_fd_sc_hd__o22a_2 _22028_ (.A1(_07560_),
    .A2(_07561_),
    .B1(_07472_),
    .B2(_07562_),
    .X(_07706_));
 sky130_fd_sc_hd__a2bb2o_2 _22029_ (.A1_N(_07705_),
    .A2_N(_07706_),
    .B1(_07705_),
    .B2(_07706_),
    .X(_07707_));
 sky130_fd_sc_hd__a2bb2o_2 _22030_ (.A1_N(_07576_),
    .A2_N(_07707_),
    .B1(_07576_),
    .B2(_07707_),
    .X(_07708_));
 sky130_fd_sc_hd__o22a_2 _22031_ (.A1(_07563_),
    .A2(_07564_),
    .B1(_07432_),
    .B2(_07565_),
    .X(_07709_));
 sky130_fd_sc_hd__a2bb2o_2 _22032_ (.A1_N(_07708_),
    .A2_N(_07709_),
    .B1(_07708_),
    .B2(_07709_),
    .X(_07710_));
 sky130_fd_sc_hd__a2bb2o_2 _22033_ (.A1_N(_07431_),
    .A2_N(_07710_),
    .B1(_07431_),
    .B2(_07710_),
    .X(_07711_));
 sky130_fd_sc_hd__o22a_2 _22034_ (.A1(_07566_),
    .A2(_07567_),
    .B1(_07428_),
    .B2(_07568_),
    .X(_07712_));
 sky130_fd_sc_hd__or2_2 _22035_ (.A(_07711_),
    .B(_07712_),
    .X(_07713_));
 sky130_vsdinv _22036_ (.A(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__a21o_2 _22037_ (.A1(_07711_),
    .A2(_07712_),
    .B1(_07714_),
    .X(_07715_));
 sky130_fd_sc_hd__a22o_2 _22038_ (.A1(_07569_),
    .A2(_07570_),
    .B1(_07418_),
    .B2(_07571_),
    .X(_07716_));
 sky130_fd_sc_hd__o31a_2 _22039_ (.A1(_07419_),
    .A2(_07572_),
    .A3(_07426_),
    .B1(_07716_),
    .X(_07717_));
 sky130_fd_sc_hd__a2bb2oi_2 _22040_ (.A1_N(_07715_),
    .A2_N(_07717_),
    .B1(_07715_),
    .B2(_07717_),
    .Y(_02653_));
 sky130_fd_sc_hd__o22a_2 _22041_ (.A1(_07708_),
    .A2(_07709_),
    .B1(_07431_),
    .B2(_07710_),
    .X(_07718_));
 sky130_vsdinv _22042_ (.A(_07718_),
    .Y(_07719_));
 sky130_fd_sc_hd__o22a_2 _22043_ (.A1(_07578_),
    .A2(_07614_),
    .B1(_07577_),
    .B2(_07615_),
    .X(_07720_));
 sky130_fd_sc_hd__o22a_2 _22044_ (.A1(_07594_),
    .A2(_07595_),
    .B1(_07579_),
    .B2(_07596_),
    .X(_07721_));
 sky130_fd_sc_hd__or2_2 _22045_ (.A(_07720_),
    .B(_07721_),
    .X(_07722_));
 sky130_fd_sc_hd__a21bo_2 _22046_ (.A1(_07720_),
    .A2(_07721_),
    .B1_N(_07722_),
    .X(_07723_));
 sky130_fd_sc_hd__o22a_2 _22047_ (.A1(_07611_),
    .A2(_07612_),
    .B1(_07597_),
    .B2(_07613_),
    .X(_07724_));
 sky130_fd_sc_hd__o22a_2 _22048_ (.A1(_07618_),
    .A2(_07645_),
    .B1(_07617_),
    .B2(_07646_),
    .X(_07725_));
 sky130_fd_sc_hd__a21oi_2 _22049_ (.A1(_07582_),
    .A2(_07584_),
    .B1(_07581_),
    .Y(_07726_));
 sky130_fd_sc_hd__buf_1 _22050_ (.A(_10585_),
    .X(_07727_));
 sky130_fd_sc_hd__buf_1 _22051_ (.A(_07727_),
    .X(_07728_));
 sky130_fd_sc_hd__nor2_2 _22052_ (.A(_07728_),
    .B(_04730_),
    .Y(_07729_));
 sky130_fd_sc_hd__a2bb2o_2 _22053_ (.A1_N(_07582_),
    .A2_N(_07729_),
    .B1(_07582_),
    .B2(_07729_),
    .X(_07730_));
 sky130_fd_sc_hd__buf_1 _22054_ (.A(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__buf_1 _22055_ (.A(_07158_),
    .X(_07732_));
 sky130_fd_sc_hd__o22a_2 _22056_ (.A1(_05171_),
    .A2(_07022_),
    .B1(_05173_),
    .B2(_07732_),
    .X(_07733_));
 sky130_fd_sc_hd__and4_2 _22057_ (.A(_05513_),
    .B(_11876_),
    .C(_05515_),
    .D(\pcpi_mul.rs1[31] ),
    .X(_07734_));
 sky130_fd_sc_hd__or2_2 _22058_ (.A(_07733_),
    .B(_07734_),
    .X(_07735_));
 sky130_vsdinv _22059_ (.A(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__a22o_2 _22060_ (.A1(_07447_),
    .A2(_07736_),
    .B1(_07295_),
    .B2(_07735_),
    .X(_07737_));
 sky130_fd_sc_hd__a21oi_2 _22061_ (.A1(_07447_),
    .A2(_07590_),
    .B1(_07588_),
    .Y(_07738_));
 sky130_fd_sc_hd__a2bb2o_2 _22062_ (.A1_N(_07737_),
    .A2_N(_07738_),
    .B1(_07737_),
    .B2(_07738_),
    .X(_07739_));
 sky130_fd_sc_hd__a2bb2o_2 _22063_ (.A1_N(_07731_),
    .A2_N(_07739_),
    .B1(_07731_),
    .B2(_07739_),
    .X(_07740_));
 sky130_fd_sc_hd__o22a_2 _22064_ (.A1(_07591_),
    .A2(_07592_),
    .B1(_07585_),
    .B2(_07593_),
    .X(_07741_));
 sky130_fd_sc_hd__a2bb2o_2 _22065_ (.A1_N(_07740_),
    .A2_N(_07741_),
    .B1(_07740_),
    .B2(_07741_),
    .X(_07742_));
 sky130_fd_sc_hd__a2bb2o_2 _22066_ (.A1_N(_07726_),
    .A2_N(_07742_),
    .B1(_07726_),
    .B2(_07742_),
    .X(_07743_));
 sky130_fd_sc_hd__o22a_2 _22067_ (.A1(_07601_),
    .A2(_07607_),
    .B1(_07600_),
    .B2(_07608_),
    .X(_07744_));
 sky130_fd_sc_hd__o22a_2 _22068_ (.A1(_07630_),
    .A2(_07631_),
    .B1(_07623_),
    .B2(_07632_),
    .X(_07745_));
 sky130_fd_sc_hd__a21oi_2 _22069_ (.A1(_07605_),
    .A2(_07606_),
    .B1(_07604_),
    .Y(_07746_));
 sky130_fd_sc_hd__o21ba_2 _22070_ (.A1(_07619_),
    .A2(_07622_),
    .B1_N(_07621_),
    .X(_07747_));
 sky130_fd_sc_hd__o22a_2 _22071_ (.A1(_07602_),
    .A2(_06624_),
    .B1(_04828_),
    .B2(_07007_),
    .X(_07748_));
 sky130_fd_sc_hd__buf_1 _22072_ (.A(\pcpi_mul.rs1[28] ),
    .X(_07749_));
 sky130_fd_sc_hd__and4_2 _22073_ (.A(_11620_),
    .B(_11884_),
    .C(_11624_),
    .D(_07749_),
    .X(_07750_));
 sky130_fd_sc_hd__nor2_2 _22074_ (.A(_07748_),
    .B(_07750_),
    .Y(_07751_));
 sky130_fd_sc_hd__nor2_2 _22075_ (.A(_04795_),
    .B(_06891_),
    .Y(_07752_));
 sky130_fd_sc_hd__a2bb2o_2 _22076_ (.A1_N(_07751_),
    .A2_N(_07752_),
    .B1(_07751_),
    .B2(_07752_),
    .X(_07753_));
 sky130_fd_sc_hd__a2bb2o_2 _22077_ (.A1_N(_07747_),
    .A2_N(_07753_),
    .B1(_07747_),
    .B2(_07753_),
    .X(_07754_));
 sky130_fd_sc_hd__a2bb2o_2 _22078_ (.A1_N(_07746_),
    .A2_N(_07754_),
    .B1(_07746_),
    .B2(_07754_),
    .X(_07755_));
 sky130_fd_sc_hd__a2bb2o_2 _22079_ (.A1_N(_07745_),
    .A2_N(_07755_),
    .B1(_07745_),
    .B2(_07755_),
    .X(_07756_));
 sky130_fd_sc_hd__a2bb2o_2 _22080_ (.A1_N(_07744_),
    .A2_N(_07756_),
    .B1(_07744_),
    .B2(_07756_),
    .X(_07757_));
 sky130_fd_sc_hd__o22a_2 _22081_ (.A1(_07599_),
    .A2(_07609_),
    .B1(_07598_),
    .B2(_07610_),
    .X(_07758_));
 sky130_fd_sc_hd__a2bb2o_2 _22082_ (.A1_N(_07757_),
    .A2_N(_07758_),
    .B1(_07757_),
    .B2(_07758_),
    .X(_07759_));
 sky130_fd_sc_hd__a2bb2o_2 _22083_ (.A1_N(_07743_),
    .A2_N(_07759_),
    .B1(_07743_),
    .B2(_07759_),
    .X(_07760_));
 sky130_fd_sc_hd__a2bb2o_2 _22084_ (.A1_N(_07725_),
    .A2_N(_07760_),
    .B1(_07725_),
    .B2(_07760_),
    .X(_07761_));
 sky130_fd_sc_hd__a2bb2o_2 _22085_ (.A1_N(_07724_),
    .A2_N(_07761_),
    .B1(_07724_),
    .B2(_07761_),
    .X(_07762_));
 sky130_fd_sc_hd__o22a_2 _22086_ (.A1(_07642_),
    .A2(_07643_),
    .B1(_07633_),
    .B2(_07644_),
    .X(_07763_));
 sky130_fd_sc_hd__o22a_2 _22087_ (.A1(_07649_),
    .A2(_07665_),
    .B1(_07648_),
    .B2(_07666_),
    .X(_07764_));
 sky130_fd_sc_hd__or2_2 _22088_ (.A(_06049_),
    .B(_06743_),
    .X(_07765_));
 sky130_fd_sc_hd__o22a_2 _22089_ (.A1(_06051_),
    .A2(_07173_),
    .B1(_06052_),
    .B2(_06376_),
    .X(_07766_));
 sky130_fd_sc_hd__and4_2 _22090_ (.A(_06054_),
    .B(_07175_),
    .C(_06055_),
    .D(_11892_),
    .X(_07767_));
 sky130_fd_sc_hd__or2_2 _22091_ (.A(_07766_),
    .B(_07767_),
    .X(_07768_));
 sky130_fd_sc_hd__a2bb2o_2 _22092_ (.A1_N(_07765_),
    .A2_N(_07768_),
    .B1(_07765_),
    .B2(_07768_),
    .X(_07769_));
 sky130_fd_sc_hd__or2_2 _22093_ (.A(_06305_),
    .B(_06359_),
    .X(_07770_));
 sky130_fd_sc_hd__o22a_2 _22094_ (.A1(_06178_),
    .A2(_05986_),
    .B1(_07481_),
    .B2(_05995_),
    .X(_07771_));
 sky130_fd_sc_hd__and4_2 _22095_ (.A(_07483_),
    .B(_06371_),
    .C(_07484_),
    .D(_11899_),
    .X(_07772_));
 sky130_fd_sc_hd__or2_2 _22096_ (.A(_07771_),
    .B(_07772_),
    .X(_07773_));
 sky130_fd_sc_hd__a2bb2o_2 _22097_ (.A1_N(_07770_),
    .A2_N(_07773_),
    .B1(_07770_),
    .B2(_07773_),
    .X(_07774_));
 sky130_fd_sc_hd__o21ba_2 _22098_ (.A1(_07625_),
    .A2(_07629_),
    .B1_N(_07628_),
    .X(_07775_));
 sky130_fd_sc_hd__a2bb2o_2 _22099_ (.A1_N(_07774_),
    .A2_N(_07775_),
    .B1(_07774_),
    .B2(_07775_),
    .X(_07776_));
 sky130_fd_sc_hd__a2bb2o_2 _22100_ (.A1_N(_07769_),
    .A2_N(_07776_),
    .B1(_07769_),
    .B2(_07776_),
    .X(_07777_));
 sky130_fd_sc_hd__o21ba_2 _22101_ (.A1(_07636_),
    .A2(_07639_),
    .B1_N(_07638_),
    .X(_07778_));
 sky130_fd_sc_hd__o21ba_2 _22102_ (.A1(_07650_),
    .A2(_07654_),
    .B1_N(_07653_),
    .X(_07779_));
 sky130_fd_sc_hd__or2_2 _22103_ (.A(_07346_),
    .B(_06237_),
    .X(_07780_));
 sky130_fd_sc_hd__o22a_2 _22104_ (.A1(_07340_),
    .A2(_06254_),
    .B1(_05392_),
    .B2(_05715_),
    .X(_07781_));
 sky130_fd_sc_hd__and4_2 _22105_ (.A(_07342_),
    .B(_06393_),
    .C(_07343_),
    .D(_11908_),
    .X(_07782_));
 sky130_fd_sc_hd__or2_2 _22106_ (.A(_07781_),
    .B(_07782_),
    .X(_07783_));
 sky130_fd_sc_hd__a2bb2o_2 _22107_ (.A1_N(_07780_),
    .A2_N(_07783_),
    .B1(_07780_),
    .B2(_07783_),
    .X(_07784_));
 sky130_fd_sc_hd__a2bb2o_2 _22108_ (.A1_N(_07779_),
    .A2_N(_07784_),
    .B1(_07779_),
    .B2(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__a2bb2o_2 _22109_ (.A1_N(_07778_),
    .A2_N(_07785_),
    .B1(_07778_),
    .B2(_07785_),
    .X(_07786_));
 sky130_fd_sc_hd__o22a_2 _22110_ (.A1(_07635_),
    .A2(_07640_),
    .B1(_07634_),
    .B2(_07641_),
    .X(_07787_));
 sky130_fd_sc_hd__a2bb2o_2 _22111_ (.A1_N(_07786_),
    .A2_N(_07787_),
    .B1(_07786_),
    .B2(_07787_),
    .X(_07788_));
 sky130_fd_sc_hd__a2bb2o_2 _22112_ (.A1_N(_07777_),
    .A2_N(_07788_),
    .B1(_07777_),
    .B2(_07788_),
    .X(_07789_));
 sky130_fd_sc_hd__a2bb2o_2 _22113_ (.A1_N(_07764_),
    .A2_N(_07789_),
    .B1(_07764_),
    .B2(_07789_),
    .X(_07790_));
 sky130_fd_sc_hd__a2bb2o_2 _22114_ (.A1_N(_07763_),
    .A2_N(_07790_),
    .B1(_07763_),
    .B2(_07790_),
    .X(_07791_));
 sky130_fd_sc_hd__o22a_2 _22115_ (.A1(_07662_),
    .A2(_07663_),
    .B1(_07655_),
    .B2(_07664_),
    .X(_07792_));
 sky130_fd_sc_hd__o22a_2 _22116_ (.A1(_07669_),
    .A2(_07675_),
    .B1(_07668_),
    .B2(_07676_),
    .X(_07793_));
 sky130_fd_sc_hd__or2_2 _22117_ (.A(_05562_),
    .B(_05510_),
    .X(_07794_));
 sky130_fd_sc_hd__o22a_2 _22118_ (.A1(_07651_),
    .A2(_05420_),
    .B1(_05659_),
    .B2(_06134_),
    .X(_07795_));
 sky130_fd_sc_hd__and4_2 _22119_ (.A(_11593_),
    .B(_05830_),
    .C(_11598_),
    .D(_06138_),
    .X(_07796_));
 sky130_fd_sc_hd__or2_2 _22120_ (.A(_07795_),
    .B(_07796_),
    .X(_07797_));
 sky130_fd_sc_hd__a2bb2o_2 _22121_ (.A1_N(_07794_),
    .A2_N(_07797_),
    .B1(_07794_),
    .B2(_07797_),
    .X(_07798_));
 sky130_fd_sc_hd__or2_2 _22122_ (.A(_07656_),
    .B(_05335_),
    .X(_07799_));
 sky130_fd_sc_hd__o22a_2 _22123_ (.A1(_07658_),
    .A2(_05740_),
    .B1(_06034_),
    .B2(_05169_),
    .X(_07800_));
 sky130_fd_sc_hd__buf_1 _22124_ (.A(_11584_),
    .X(_07801_));
 sky130_fd_sc_hd__buf_1 _22125_ (.A(_11588_),
    .X(_07802_));
 sky130_fd_sc_hd__and4_2 _22126_ (.A(_07801_),
    .B(_11925_),
    .C(_07802_),
    .D(_05848_),
    .X(_07803_));
 sky130_fd_sc_hd__or2_2 _22127_ (.A(_07800_),
    .B(_07803_),
    .X(_07804_));
 sky130_fd_sc_hd__a2bb2o_2 _22128_ (.A1_N(_07799_),
    .A2_N(_07804_),
    .B1(_07799_),
    .B2(_07804_),
    .X(_07805_));
 sky130_fd_sc_hd__o21ba_2 _22129_ (.A1(_07657_),
    .A2(_07661_),
    .B1_N(_07660_),
    .X(_07806_));
 sky130_fd_sc_hd__a2bb2o_2 _22130_ (.A1_N(_07805_),
    .A2_N(_07806_),
    .B1(_07805_),
    .B2(_07806_),
    .X(_07807_));
 sky130_fd_sc_hd__a2bb2o_2 _22131_ (.A1_N(_07798_),
    .A2_N(_07807_),
    .B1(_07798_),
    .B2(_07807_),
    .X(_07808_));
 sky130_fd_sc_hd__a2bb2o_2 _22132_ (.A1_N(_07793_),
    .A2_N(_07808_),
    .B1(_07793_),
    .B2(_07808_),
    .X(_07809_));
 sky130_fd_sc_hd__a2bb2o_2 _22133_ (.A1_N(_07792_),
    .A2_N(_07809_),
    .B1(_07792_),
    .B2(_07809_),
    .X(_07810_));
 sky130_fd_sc_hd__o21ba_2 _22134_ (.A1(_07670_),
    .A2(_07674_),
    .B1_N(_07673_),
    .X(_07811_));
 sky130_fd_sc_hd__o21ba_2 _22135_ (.A1(_07678_),
    .A2(_07683_),
    .B1_N(_07682_),
    .X(_07812_));
 sky130_fd_sc_hd__or2_2 _22136_ (.A(_06447_),
    .B(_05155_),
    .X(_07813_));
 sky130_fd_sc_hd__buf_1 _22137_ (.A(_06974_),
    .X(_07814_));
 sky130_fd_sc_hd__o22a_2 _22138_ (.A1(_07814_),
    .A2(_05943_),
    .B1(_06445_),
    .B2(_05070_),
    .X(_07815_));
 sky130_fd_sc_hd__buf_1 _22139_ (.A(_11574_),
    .X(_07816_));
 sky130_fd_sc_hd__and4_2 _22140_ (.A(_07816_),
    .B(_11931_),
    .C(_07672_),
    .D(_11929_),
    .X(_07817_));
 sky130_fd_sc_hd__or2_2 _22141_ (.A(_07815_),
    .B(_07817_),
    .X(_07818_));
 sky130_fd_sc_hd__a2bb2o_2 _22142_ (.A1_N(_07813_),
    .A2_N(_07818_),
    .B1(_07813_),
    .B2(_07818_),
    .X(_07819_));
 sky130_fd_sc_hd__a2bb2o_2 _22143_ (.A1_N(_07812_),
    .A2_N(_07819_),
    .B1(_07812_),
    .B2(_07819_),
    .X(_07820_));
 sky130_fd_sc_hd__a2bb2o_2 _22144_ (.A1_N(_07811_),
    .A2_N(_07820_),
    .B1(_07811_),
    .B2(_07820_),
    .X(_07821_));
 sky130_fd_sc_hd__buf_1 _22145_ (.A(_06685_),
    .X(_07822_));
 sky130_fd_sc_hd__or2_2 _22146_ (.A(_07822_),
    .B(_06568_),
    .X(_07823_));
 sky130_fd_sc_hd__o22a_2 _22147_ (.A1(_07535_),
    .A2(_06277_),
    .B1(_07536_),
    .B2(_05396_),
    .X(_07824_));
 sky130_fd_sc_hd__and4_2 _22148_ (.A(_07538_),
    .B(_11940_),
    .C(_07681_),
    .D(_11937_),
    .X(_07825_));
 sky130_fd_sc_hd__or2_2 _22149_ (.A(_07824_),
    .B(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__a2bb2o_2 _22150_ (.A1_N(_07823_),
    .A2_N(_07826_),
    .B1(_07823_),
    .B2(_07826_),
    .X(_07827_));
 sky130_fd_sc_hd__buf_1 _22151_ (.A(_07099_),
    .X(_07828_));
 sky130_fd_sc_hd__or2_2 _22152_ (.A(_07828_),
    .B(_06151_),
    .X(_07829_));
 sky130_fd_sc_hd__buf_1 _22153_ (.A(_07393_),
    .X(_07830_));
 sky130_fd_sc_hd__and4_2 _22154_ (.A(_07830_),
    .B(_05406_),
    .C(_11560_),
    .D(_11946_),
    .X(_07831_));
 sky130_fd_sc_hd__buf_1 _22155_ (.A(_10596_),
    .X(_07832_));
 sky130_fd_sc_hd__o22a_2 _22156_ (.A1(_07832_),
    .A2(_11949_),
    .B1(_07247_),
    .B2(_05137_),
    .X(_07833_));
 sky130_fd_sc_hd__or2_2 _22157_ (.A(_07831_),
    .B(_07833_),
    .X(_07834_));
 sky130_fd_sc_hd__a2bb2o_2 _22158_ (.A1_N(_07829_),
    .A2_N(_07834_),
    .B1(_07829_),
    .B2(_07834_),
    .X(_07835_));
 sky130_fd_sc_hd__o21ba_2 _22159_ (.A1(_07685_),
    .A2(_07689_),
    .B1_N(_07687_),
    .X(_07836_));
 sky130_fd_sc_hd__a2bb2o_2 _22160_ (.A1_N(_07835_),
    .A2_N(_07836_),
    .B1(_07835_),
    .B2(_07836_),
    .X(_07837_));
 sky130_fd_sc_hd__a2bb2o_2 _22161_ (.A1_N(_07827_),
    .A2_N(_07837_),
    .B1(_07827_),
    .B2(_07837_),
    .X(_07838_));
 sky130_fd_sc_hd__o22a_2 _22162_ (.A1(_07690_),
    .A2(_07691_),
    .B1(_07684_),
    .B2(_07692_),
    .X(_07839_));
 sky130_fd_sc_hd__a2bb2o_2 _22163_ (.A1_N(_07838_),
    .A2_N(_07839_),
    .B1(_07838_),
    .B2(_07839_),
    .X(_07840_));
 sky130_fd_sc_hd__a2bb2o_2 _22164_ (.A1_N(_07821_),
    .A2_N(_07840_),
    .B1(_07821_),
    .B2(_07840_),
    .X(_07841_));
 sky130_fd_sc_hd__o22a_2 _22165_ (.A1(_07693_),
    .A2(_07694_),
    .B1(_07677_),
    .B2(_07695_),
    .X(_07842_));
 sky130_fd_sc_hd__a2bb2o_2 _22166_ (.A1_N(_07841_),
    .A2_N(_07842_),
    .B1(_07841_),
    .B2(_07842_),
    .X(_07843_));
 sky130_fd_sc_hd__a2bb2o_2 _22167_ (.A1_N(_07810_),
    .A2_N(_07843_),
    .B1(_07810_),
    .B2(_07843_),
    .X(_07844_));
 sky130_fd_sc_hd__o22a_2 _22168_ (.A1(_07696_),
    .A2(_07697_),
    .B1(_07667_),
    .B2(_07698_),
    .X(_07845_));
 sky130_fd_sc_hd__a2bb2o_2 _22169_ (.A1_N(_07844_),
    .A2_N(_07845_),
    .B1(_07844_),
    .B2(_07845_),
    .X(_07846_));
 sky130_fd_sc_hd__a2bb2o_2 _22170_ (.A1_N(_07791_),
    .A2_N(_07846_),
    .B1(_07791_),
    .B2(_07846_),
    .X(_07847_));
 sky130_fd_sc_hd__o22a_2 _22171_ (.A1(_07699_),
    .A2(_07700_),
    .B1(_07647_),
    .B2(_07701_),
    .X(_07848_));
 sky130_fd_sc_hd__a2bb2o_2 _22172_ (.A1_N(_07847_),
    .A2_N(_07848_),
    .B1(_07847_),
    .B2(_07848_),
    .X(_07849_));
 sky130_fd_sc_hd__a2bb2o_2 _22173_ (.A1_N(_07762_),
    .A2_N(_07849_),
    .B1(_07762_),
    .B2(_07849_),
    .X(_07850_));
 sky130_fd_sc_hd__o22a_2 _22174_ (.A1(_07702_),
    .A2(_07703_),
    .B1(_07616_),
    .B2(_07704_),
    .X(_07851_));
 sky130_fd_sc_hd__a2bb2o_2 _22175_ (.A1_N(_07850_),
    .A2_N(_07851_),
    .B1(_07850_),
    .B2(_07851_),
    .X(_07852_));
 sky130_fd_sc_hd__a2bb2o_2 _22176_ (.A1_N(_07723_),
    .A2_N(_07852_),
    .B1(_07723_),
    .B2(_07852_),
    .X(_07853_));
 sky130_fd_sc_hd__o22a_2 _22177_ (.A1(_07705_),
    .A2(_07706_),
    .B1(_07576_),
    .B2(_07707_),
    .X(_07854_));
 sky130_fd_sc_hd__a2bb2o_2 _22178_ (.A1_N(_07853_),
    .A2_N(_07854_),
    .B1(_07853_),
    .B2(_07854_),
    .X(_07855_));
 sky130_fd_sc_hd__a2bb2o_2 _22179_ (.A1_N(_07575_),
    .A2_N(_07855_),
    .B1(_07575_),
    .B2(_07855_),
    .X(_07856_));
 sky130_vsdinv _22180_ (.A(_07856_),
    .Y(_07857_));
 sky130_fd_sc_hd__a22o_2 _22181_ (.A1(_07719_),
    .A2(_07857_),
    .B1(_07718_),
    .B2(_07856_),
    .X(_07858_));
 sky130_fd_sc_hd__o21ai_2 _22182_ (.A1(_07715_),
    .A2(_07717_),
    .B1(_07713_),
    .Y(_07859_));
 sky130_fd_sc_hd__a2bb2o_2 _22183_ (.A1_N(_07858_),
    .A2_N(_07859_),
    .B1(_07858_),
    .B2(_07859_),
    .X(_02654_));
 sky130_fd_sc_hd__o22a_2 _22184_ (.A1(_07725_),
    .A2(_07760_),
    .B1(_07724_),
    .B2(_07761_),
    .X(_07860_));
 sky130_fd_sc_hd__o22a_2 _22185_ (.A1(_07740_),
    .A2(_07741_),
    .B1(_07726_),
    .B2(_07742_),
    .X(_07861_));
 sky130_fd_sc_hd__or2_2 _22186_ (.A(_07860_),
    .B(_07861_),
    .X(_07862_));
 sky130_fd_sc_hd__a21bo_2 _22187_ (.A1(_07860_),
    .A2(_07861_),
    .B1_N(_07862_),
    .X(_07863_));
 sky130_fd_sc_hd__o22a_2 _22188_ (.A1(_07757_),
    .A2(_07758_),
    .B1(_07743_),
    .B2(_07759_),
    .X(_07864_));
 sky130_fd_sc_hd__o22a_2 _22189_ (.A1(_07764_),
    .A2(_07789_),
    .B1(_07763_),
    .B2(_07790_),
    .X(_07865_));
 sky130_fd_sc_hd__a21oi_2 _22190_ (.A1(_07582_),
    .A2(_07729_),
    .B1(_07581_),
    .Y(_07866_));
 sky130_fd_sc_hd__buf_1 _22191_ (.A(_07866_),
    .X(_07867_));
 sky130_fd_sc_hd__buf_1 _22192_ (.A(\pcpi_mul.rs1[32] ),
    .X(_07868_));
 sky130_fd_sc_hd__buf_1 _22193_ (.A(_07868_),
    .X(_07869_));
 sky130_fd_sc_hd__buf_1 _22194_ (.A(_07869_),
    .X(_07870_));
 sky130_fd_sc_hd__a31o_2 _22195_ (.A1(_07870_),
    .A2(\pcpi_mul.rs2[0] ),
    .A3(_07736_),
    .B1(_07734_),
    .X(_07871_));
 sky130_vsdinv _22196_ (.A(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__o22a_2 _22197_ (.A1(_06368_),
    .A2(_07159_),
    .B1(_10586_),
    .B2(_06369_),
    .X(_07873_));
 sky130_fd_sc_hd__and4_2 _22198_ (.A(_06115_),
    .B(_11873_),
    .C(_07868_),
    .D(_06116_),
    .X(_07874_));
 sky130_fd_sc_hd__nor2_2 _22199_ (.A(_07873_),
    .B(_07874_),
    .Y(_07875_));
 sky130_fd_sc_hd__o2bb2a_2 _22200_ (.A1_N(_07297_),
    .A2_N(_07875_),
    .B1(_07297_),
    .B2(_07875_),
    .X(_07876_));
 sky130_vsdinv _22201_ (.A(_07876_),
    .Y(_07877_));
 sky130_fd_sc_hd__a22o_2 _22202_ (.A1(_07872_),
    .A2(_07877_),
    .B1(_07871_),
    .B2(_07876_),
    .X(_07878_));
 sky130_fd_sc_hd__a2bb2o_2 _22203_ (.A1_N(_07730_),
    .A2_N(_07878_),
    .B1(_07730_),
    .B2(_07878_),
    .X(_07879_));
 sky130_fd_sc_hd__o22a_2 _22204_ (.A1(_07737_),
    .A2(_07738_),
    .B1(_07730_),
    .B2(_07739_),
    .X(_07880_));
 sky130_fd_sc_hd__a2bb2o_2 _22205_ (.A1_N(_07879_),
    .A2_N(_07880_),
    .B1(_07879_),
    .B2(_07880_),
    .X(_07881_));
 sky130_fd_sc_hd__a2bb2o_2 _22206_ (.A1_N(_07867_),
    .A2_N(_07881_),
    .B1(_07867_),
    .B2(_07881_),
    .X(_07882_));
 sky130_fd_sc_hd__o22a_2 _22207_ (.A1(_07747_),
    .A2(_07753_),
    .B1(_07746_),
    .B2(_07754_),
    .X(_07883_));
 sky130_fd_sc_hd__o22a_2 _22208_ (.A1(_07774_),
    .A2(_07775_),
    .B1(_07769_),
    .B2(_07776_),
    .X(_07884_));
 sky130_fd_sc_hd__a21oi_2 _22209_ (.A1(_07751_),
    .A2(_07752_),
    .B1(_07750_),
    .Y(_07885_));
 sky130_fd_sc_hd__o21ba_2 _22210_ (.A1(_07765_),
    .A2(_07768_),
    .B1_N(_07767_),
    .X(_07886_));
 sky130_fd_sc_hd__o22a_2 _22211_ (.A1(_07602_),
    .A2(_06749_),
    .B1(_04828_),
    .B2(_07009_),
    .X(_07887_));
 sky130_fd_sc_hd__and4_2 _22212_ (.A(_11620_),
    .B(_07749_),
    .C(_11624_),
    .D(_07587_),
    .X(_07888_));
 sky130_fd_sc_hd__nor2_2 _22213_ (.A(_07887_),
    .B(_07888_),
    .Y(_07889_));
 sky130_fd_sc_hd__nor2_2 _22214_ (.A(_04795_),
    .B(_07285_),
    .Y(_07890_));
 sky130_fd_sc_hd__a2bb2o_2 _22215_ (.A1_N(_07889_),
    .A2_N(_07890_),
    .B1(_07889_),
    .B2(_07890_),
    .X(_07891_));
 sky130_fd_sc_hd__a2bb2o_2 _22216_ (.A1_N(_07886_),
    .A2_N(_07891_),
    .B1(_07886_),
    .B2(_07891_),
    .X(_07892_));
 sky130_fd_sc_hd__a2bb2o_2 _22217_ (.A1_N(_07885_),
    .A2_N(_07892_),
    .B1(_07885_),
    .B2(_07892_),
    .X(_07893_));
 sky130_fd_sc_hd__a2bb2o_2 _22218_ (.A1_N(_07884_),
    .A2_N(_07893_),
    .B1(_07884_),
    .B2(_07893_),
    .X(_07894_));
 sky130_fd_sc_hd__a2bb2o_2 _22219_ (.A1_N(_07883_),
    .A2_N(_07894_),
    .B1(_07883_),
    .B2(_07894_),
    .X(_07895_));
 sky130_fd_sc_hd__o22a_2 _22220_ (.A1(_07745_),
    .A2(_07755_),
    .B1(_07744_),
    .B2(_07756_),
    .X(_07896_));
 sky130_fd_sc_hd__a2bb2o_2 _22221_ (.A1_N(_07895_),
    .A2_N(_07896_),
    .B1(_07895_),
    .B2(_07896_),
    .X(_07897_));
 sky130_fd_sc_hd__a2bb2o_2 _22222_ (.A1_N(_07882_),
    .A2_N(_07897_),
    .B1(_07882_),
    .B2(_07897_),
    .X(_07898_));
 sky130_fd_sc_hd__a2bb2o_2 _22223_ (.A1_N(_07865_),
    .A2_N(_07898_),
    .B1(_07865_),
    .B2(_07898_),
    .X(_07899_));
 sky130_fd_sc_hd__a2bb2o_2 _22224_ (.A1_N(_07864_),
    .A2_N(_07899_),
    .B1(_07864_),
    .B2(_07899_),
    .X(_07900_));
 sky130_fd_sc_hd__o22a_2 _22225_ (.A1(_07786_),
    .A2(_07787_),
    .B1(_07777_),
    .B2(_07788_),
    .X(_07901_));
 sky130_fd_sc_hd__o22a_2 _22226_ (.A1(_07793_),
    .A2(_07808_),
    .B1(_07792_),
    .B2(_07809_),
    .X(_07902_));
 sky130_fd_sc_hd__or2_2 _22227_ (.A(_06049_),
    .B(_06879_),
    .X(_07903_));
 sky130_fd_sc_hd__o22a_2 _22228_ (.A1(_06051_),
    .A2(_06376_),
    .B1(_04951_),
    .B2(_06742_),
    .X(_07904_));
 sky130_fd_sc_hd__and4_2 _22229_ (.A(_11614_),
    .B(_11892_),
    .C(_11617_),
    .D(_07459_),
    .X(_07905_));
 sky130_fd_sc_hd__or2_2 _22230_ (.A(_07904_),
    .B(_07905_),
    .X(_07906_));
 sky130_fd_sc_hd__a2bb2o_2 _22231_ (.A1_N(_07903_),
    .A2_N(_07906_),
    .B1(_07903_),
    .B2(_07906_),
    .X(_07907_));
 sky130_fd_sc_hd__or2_2 _22232_ (.A(_07624_),
    .B(_06361_),
    .X(_07908_));
 sky130_fd_sc_hd__o22a_2 _22233_ (.A1(_07626_),
    .A2(_05995_),
    .B1(_05132_),
    .B2(_06111_),
    .X(_07909_));
 sky130_fd_sc_hd__and4_2 _22234_ (.A(_11608_),
    .B(_11899_),
    .C(_11611_),
    .D(_07038_),
    .X(_07910_));
 sky130_fd_sc_hd__or2_2 _22235_ (.A(_07909_),
    .B(_07910_),
    .X(_07911_));
 sky130_fd_sc_hd__a2bb2o_2 _22236_ (.A1_N(_07908_),
    .A2_N(_07911_),
    .B1(_07908_),
    .B2(_07911_),
    .X(_07912_));
 sky130_fd_sc_hd__o21ba_2 _22237_ (.A1(_07770_),
    .A2(_07773_),
    .B1_N(_07772_),
    .X(_07913_));
 sky130_fd_sc_hd__a2bb2o_2 _22238_ (.A1_N(_07912_),
    .A2_N(_07913_),
    .B1(_07912_),
    .B2(_07913_),
    .X(_07914_));
 sky130_fd_sc_hd__a2bb2o_2 _22239_ (.A1_N(_07907_),
    .A2_N(_07914_),
    .B1(_07907_),
    .B2(_07914_),
    .X(_07915_));
 sky130_fd_sc_hd__o21ba_2 _22240_ (.A1(_07780_),
    .A2(_07783_),
    .B1_N(_07782_),
    .X(_07916_));
 sky130_fd_sc_hd__o21ba_2 _22241_ (.A1(_07794_),
    .A2(_07797_),
    .B1_N(_07796_),
    .X(_07917_));
 sky130_fd_sc_hd__buf_1 _22242_ (.A(_06318_),
    .X(_07918_));
 sky130_fd_sc_hd__o22a_2 _22243_ (.A1(_07918_),
    .A2(_07196_),
    .B1(_05389_),
    .B2(_05884_),
    .X(_07919_));
 sky130_fd_sc_hd__and4_2 _22244_ (.A(_11603_),
    .B(_06117_),
    .C(_11606_),
    .D(_11905_),
    .X(_07920_));
 sky130_fd_sc_hd__nor2_2 _22245_ (.A(_07919_),
    .B(_07920_),
    .Y(_07921_));
 sky130_fd_sc_hd__buf_1 _22246_ (.A(_05393_),
    .X(_07922_));
 sky130_fd_sc_hd__nor2_2 _22247_ (.A(_07922_),
    .B(_05988_),
    .Y(_07923_));
 sky130_fd_sc_hd__a2bb2o_2 _22248_ (.A1_N(_07921_),
    .A2_N(_07923_),
    .B1(_07921_),
    .B2(_07923_),
    .X(_07924_));
 sky130_fd_sc_hd__a2bb2o_2 _22249_ (.A1_N(_07917_),
    .A2_N(_07924_),
    .B1(_07917_),
    .B2(_07924_),
    .X(_07925_));
 sky130_fd_sc_hd__a2bb2o_2 _22250_ (.A1_N(_07916_),
    .A2_N(_07925_),
    .B1(_07916_),
    .B2(_07925_),
    .X(_07926_));
 sky130_fd_sc_hd__o22a_2 _22251_ (.A1(_07779_),
    .A2(_07784_),
    .B1(_07778_),
    .B2(_07785_),
    .X(_07927_));
 sky130_fd_sc_hd__a2bb2o_2 _22252_ (.A1_N(_07926_),
    .A2_N(_07927_),
    .B1(_07926_),
    .B2(_07927_),
    .X(_07928_));
 sky130_fd_sc_hd__a2bb2o_2 _22253_ (.A1_N(_07915_),
    .A2_N(_07928_),
    .B1(_07915_),
    .B2(_07928_),
    .X(_07929_));
 sky130_fd_sc_hd__a2bb2o_2 _22254_ (.A1_N(_07902_),
    .A2_N(_07929_),
    .B1(_07902_),
    .B2(_07929_),
    .X(_07930_));
 sky130_fd_sc_hd__a2bb2o_2 _22255_ (.A1_N(_07901_),
    .A2_N(_07930_),
    .B1(_07901_),
    .B2(_07930_),
    .X(_07931_));
 sky130_fd_sc_hd__o22a_2 _22256_ (.A1(_07805_),
    .A2(_07806_),
    .B1(_07798_),
    .B2(_07807_),
    .X(_07932_));
 sky130_fd_sc_hd__o22a_2 _22257_ (.A1(_07812_),
    .A2(_07819_),
    .B1(_07811_),
    .B2(_07820_),
    .X(_07933_));
 sky130_fd_sc_hd__or2_2 _22258_ (.A(_05562_),
    .B(_06255_),
    .X(_07934_));
 sky130_fd_sc_hd__o22a_2 _22259_ (.A1(_07651_),
    .A2(_05501_),
    .B1(_05659_),
    .B2(_05598_),
    .X(_07935_));
 sky130_fd_sc_hd__and4_2 _22260_ (.A(_11593_),
    .B(_05831_),
    .C(_11598_),
    .D(_06392_),
    .X(_07936_));
 sky130_fd_sc_hd__or2_2 _22261_ (.A(_07935_),
    .B(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__a2bb2o_2 _22262_ (.A1_N(_07934_),
    .A2_N(_07937_),
    .B1(_07934_),
    .B2(_07937_),
    .X(_07938_));
 sky130_fd_sc_hd__or2_2 _22263_ (.A(_07656_),
    .B(_05421_),
    .X(_07939_));
 sky130_fd_sc_hd__o22a_2 _22264_ (.A1(_07658_),
    .A2(_05169_),
    .B1(_06034_),
    .B2(_05334_),
    .X(_07940_));
 sky130_fd_sc_hd__and4_2 _22265_ (.A(_07515_),
    .B(_05848_),
    .C(_07516_),
    .D(_07509_),
    .X(_07941_));
 sky130_fd_sc_hd__or2_2 _22266_ (.A(_07940_),
    .B(_07941_),
    .X(_07942_));
 sky130_fd_sc_hd__a2bb2o_2 _22267_ (.A1_N(_07939_),
    .A2_N(_07942_),
    .B1(_07939_),
    .B2(_07942_),
    .X(_07943_));
 sky130_fd_sc_hd__o21ba_2 _22268_ (.A1(_07799_),
    .A2(_07804_),
    .B1_N(_07803_),
    .X(_07944_));
 sky130_fd_sc_hd__a2bb2o_2 _22269_ (.A1_N(_07943_),
    .A2_N(_07944_),
    .B1(_07943_),
    .B2(_07944_),
    .X(_07945_));
 sky130_fd_sc_hd__a2bb2o_2 _22270_ (.A1_N(_07938_),
    .A2_N(_07945_),
    .B1(_07938_),
    .B2(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__a2bb2o_2 _22271_ (.A1_N(_07933_),
    .A2_N(_07946_),
    .B1(_07933_),
    .B2(_07946_),
    .X(_07947_));
 sky130_fd_sc_hd__a2bb2o_2 _22272_ (.A1_N(_07932_),
    .A2_N(_07947_),
    .B1(_07932_),
    .B2(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__o21ba_2 _22273_ (.A1(_07813_),
    .A2(_07818_),
    .B1_N(_07817_),
    .X(_07949_));
 sky130_fd_sc_hd__o21ba_2 _22274_ (.A1(_07823_),
    .A2(_07826_),
    .B1_N(_07825_),
    .X(_07950_));
 sky130_fd_sc_hd__or2_2 _22275_ (.A(_07376_),
    .B(_05158_),
    .X(_07951_));
 sky130_fd_sc_hd__o22a_2 _22276_ (.A1(_07378_),
    .A2(_05070_),
    .B1(_07379_),
    .B2(_05072_),
    .X(_07952_));
 sky130_fd_sc_hd__and4_2 _22277_ (.A(_07816_),
    .B(_11929_),
    .C(_07672_),
    .D(_11927_),
    .X(_07953_));
 sky130_fd_sc_hd__or2_2 _22278_ (.A(_07952_),
    .B(_07953_),
    .X(_07954_));
 sky130_fd_sc_hd__a2bb2o_2 _22279_ (.A1_N(_07951_),
    .A2_N(_07954_),
    .B1(_07951_),
    .B2(_07954_),
    .X(_07955_));
 sky130_fd_sc_hd__a2bb2o_2 _22280_ (.A1_N(_07950_),
    .A2_N(_07955_),
    .B1(_07950_),
    .B2(_07955_),
    .X(_07956_));
 sky130_fd_sc_hd__a2bb2o_2 _22281_ (.A1_N(_07949_),
    .A2_N(_07956_),
    .B1(_07949_),
    .B2(_07956_),
    .X(_07957_));
 sky130_fd_sc_hd__or2_2 _22282_ (.A(_06686_),
    .B(_05077_),
    .X(_07958_));
 sky130_fd_sc_hd__o22a_2 _22283_ (.A1(_07535_),
    .A2(_05396_),
    .B1(_07536_),
    .B2(_05017_),
    .X(_07959_));
 sky130_fd_sc_hd__and4_2 _22284_ (.A(_07538_),
    .B(_11937_),
    .C(_07539_),
    .D(_11934_),
    .X(_07960_));
 sky130_fd_sc_hd__or2_2 _22285_ (.A(_07959_),
    .B(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__a2bb2o_2 _22286_ (.A1_N(_07958_),
    .A2_N(_07961_),
    .B1(_07958_),
    .B2(_07961_),
    .X(_07962_));
 sky130_fd_sc_hd__or2_2 _22287_ (.A(_07828_),
    .B(_06277_),
    .X(_07963_));
 sky130_fd_sc_hd__and4_2 _22288_ (.A(_07830_),
    .B(_05137_),
    .C(_11560_),
    .D(_05197_),
    .X(_07964_));
 sky130_fd_sc_hd__buf_1 _22289_ (.A(_07246_),
    .X(_07965_));
 sky130_fd_sc_hd__o22a_2 _22290_ (.A1(_07832_),
    .A2(_11946_),
    .B1(_07965_),
    .B2(_05194_),
    .X(_07966_));
 sky130_fd_sc_hd__or2_2 _22291_ (.A(_07964_),
    .B(_07966_),
    .X(_07967_));
 sky130_fd_sc_hd__a2bb2o_2 _22292_ (.A1_N(_07963_),
    .A2_N(_07967_),
    .B1(_07963_),
    .B2(_07967_),
    .X(_07968_));
 sky130_fd_sc_hd__o21ba_2 _22293_ (.A1(_07829_),
    .A2(_07834_),
    .B1_N(_07831_),
    .X(_07969_));
 sky130_fd_sc_hd__a2bb2o_2 _22294_ (.A1_N(_07968_),
    .A2_N(_07969_),
    .B1(_07968_),
    .B2(_07969_),
    .X(_07970_));
 sky130_fd_sc_hd__a2bb2o_2 _22295_ (.A1_N(_07962_),
    .A2_N(_07970_),
    .B1(_07962_),
    .B2(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__o22a_2 _22296_ (.A1(_07835_),
    .A2(_07836_),
    .B1(_07827_),
    .B2(_07837_),
    .X(_07972_));
 sky130_fd_sc_hd__a2bb2o_2 _22297_ (.A1_N(_07971_),
    .A2_N(_07972_),
    .B1(_07971_),
    .B2(_07972_),
    .X(_07973_));
 sky130_fd_sc_hd__a2bb2o_2 _22298_ (.A1_N(_07957_),
    .A2_N(_07973_),
    .B1(_07957_),
    .B2(_07973_),
    .X(_07974_));
 sky130_fd_sc_hd__o22a_2 _22299_ (.A1(_07838_),
    .A2(_07839_),
    .B1(_07821_),
    .B2(_07840_),
    .X(_07975_));
 sky130_fd_sc_hd__a2bb2o_2 _22300_ (.A1_N(_07974_),
    .A2_N(_07975_),
    .B1(_07974_),
    .B2(_07975_),
    .X(_07976_));
 sky130_fd_sc_hd__a2bb2o_2 _22301_ (.A1_N(_07948_),
    .A2_N(_07976_),
    .B1(_07948_),
    .B2(_07976_),
    .X(_07977_));
 sky130_fd_sc_hd__o22a_2 _22302_ (.A1(_07841_),
    .A2(_07842_),
    .B1(_07810_),
    .B2(_07843_),
    .X(_07978_));
 sky130_fd_sc_hd__a2bb2o_2 _22303_ (.A1_N(_07977_),
    .A2_N(_07978_),
    .B1(_07977_),
    .B2(_07978_),
    .X(_07979_));
 sky130_fd_sc_hd__a2bb2o_2 _22304_ (.A1_N(_07931_),
    .A2_N(_07979_),
    .B1(_07931_),
    .B2(_07979_),
    .X(_07980_));
 sky130_fd_sc_hd__o22a_2 _22305_ (.A1(_07844_),
    .A2(_07845_),
    .B1(_07791_),
    .B2(_07846_),
    .X(_07981_));
 sky130_fd_sc_hd__a2bb2o_2 _22306_ (.A1_N(_07980_),
    .A2_N(_07981_),
    .B1(_07980_),
    .B2(_07981_),
    .X(_07982_));
 sky130_fd_sc_hd__a2bb2o_2 _22307_ (.A1_N(_07900_),
    .A2_N(_07982_),
    .B1(_07900_),
    .B2(_07982_),
    .X(_07983_));
 sky130_fd_sc_hd__o22a_2 _22308_ (.A1(_07847_),
    .A2(_07848_),
    .B1(_07762_),
    .B2(_07849_),
    .X(_07984_));
 sky130_fd_sc_hd__a2bb2o_2 _22309_ (.A1_N(_07983_),
    .A2_N(_07984_),
    .B1(_07983_),
    .B2(_07984_),
    .X(_07985_));
 sky130_fd_sc_hd__a2bb2o_2 _22310_ (.A1_N(_07863_),
    .A2_N(_07985_),
    .B1(_07863_),
    .B2(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__o22a_2 _22311_ (.A1(_07850_),
    .A2(_07851_),
    .B1(_07723_),
    .B2(_07852_),
    .X(_07987_));
 sky130_fd_sc_hd__a2bb2o_2 _22312_ (.A1_N(_07986_),
    .A2_N(_07987_),
    .B1(_07986_),
    .B2(_07987_),
    .X(_07988_));
 sky130_fd_sc_hd__a2bb2o_2 _22313_ (.A1_N(_07722_),
    .A2_N(_07988_),
    .B1(_07722_),
    .B2(_07988_),
    .X(_07989_));
 sky130_fd_sc_hd__o22a_2 _22314_ (.A1(_07853_),
    .A2(_07854_),
    .B1(_07575_),
    .B2(_07855_),
    .X(_07990_));
 sky130_fd_sc_hd__or2_2 _22315_ (.A(_07989_),
    .B(_07990_),
    .X(_07991_));
 sky130_fd_sc_hd__a21bo_2 _22316_ (.A1(_07989_),
    .A2(_07990_),
    .B1_N(_07991_),
    .X(_07992_));
 sky130_fd_sc_hd__or2_2 _22317_ (.A(_07715_),
    .B(_07858_),
    .X(_07993_));
 sky130_fd_sc_hd__or3_2 _22318_ (.A(_07419_),
    .B(_07572_),
    .C(_07993_),
    .X(_07994_));
 sky130_fd_sc_hd__o21ai_2 _22319_ (.A1(_07719_),
    .A2(_07857_),
    .B1(_07714_),
    .Y(_07995_));
 sky130_fd_sc_hd__o221a_2 _22320_ (.A1(_07718_),
    .A2(_07856_),
    .B1(_07716_),
    .B2(_07993_),
    .C1(_07995_),
    .X(_07996_));
 sky130_fd_sc_hd__o21ai_2 _22321_ (.A1(_07426_),
    .A2(_07994_),
    .B1(_07996_),
    .Y(_07997_));
 sky130_vsdinv _22322_ (.A(_07997_),
    .Y(_07998_));
 sky130_vsdinv _22323_ (.A(_07992_),
    .Y(_07999_));
 sky130_fd_sc_hd__o22a_2 _22324_ (.A1(_07992_),
    .A2(_07998_),
    .B1(_07999_),
    .B2(_07997_),
    .X(_02655_));
 sky130_fd_sc_hd__o22a_2 _22325_ (.A1(_07986_),
    .A2(_07987_),
    .B1(_07722_),
    .B2(_07988_),
    .X(_08000_));
 sky130_fd_sc_hd__o22a_2 _22326_ (.A1(_07865_),
    .A2(_07898_),
    .B1(_07864_),
    .B2(_07899_),
    .X(_08001_));
 sky130_fd_sc_hd__buf_1 _22327_ (.A(_07867_),
    .X(_08002_));
 sky130_fd_sc_hd__o22a_2 _22328_ (.A1(_07879_),
    .A2(_07880_),
    .B1(_08002_),
    .B2(_07881_),
    .X(_08003_));
 sky130_fd_sc_hd__or2_2 _22329_ (.A(_08001_),
    .B(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__a21bo_2 _22330_ (.A1(_08001_),
    .A2(_08003_),
    .B1_N(_08004_),
    .X(_08005_));
 sky130_fd_sc_hd__o22a_2 _22331_ (.A1(_07895_),
    .A2(_07896_),
    .B1(_07882_),
    .B2(_07897_),
    .X(_08006_));
 sky130_fd_sc_hd__o22a_2 _22332_ (.A1(_07902_),
    .A2(_07929_),
    .B1(_07901_),
    .B2(_07930_),
    .X(_08007_));
 sky130_fd_sc_hd__o22a_2 _22333_ (.A1(_07872_),
    .A2(_07877_),
    .B1(_07731_),
    .B2(_07878_),
    .X(_08008_));
 sky130_fd_sc_hd__or4_2 _22334_ (.A(_10587_),
    .B(_06369_),
    .C(_07728_),
    .D(_06368_),
    .X(_08009_));
 sky130_fd_sc_hd__a22o_2 _22335_ (.A1(_07869_),
    .A2(_11633_),
    .B1(_07869_),
    .B2(_11629_),
    .X(_08010_));
 sky130_fd_sc_hd__nand2_2 _22336_ (.A(_08009_),
    .B(_08010_),
    .Y(_08011_));
 sky130_fd_sc_hd__o22a_2 _22337_ (.A1(_07447_),
    .A2(_07874_),
    .B1(_04539_),
    .B2(_07873_),
    .X(_08012_));
 sky130_fd_sc_hd__a2bb2o_2 _22338_ (.A1_N(_08011_),
    .A2_N(_08012_),
    .B1(_08011_),
    .B2(_08012_),
    .X(_08013_));
 sky130_fd_sc_hd__nor2_2 _22339_ (.A(_07731_),
    .B(_08013_),
    .Y(_08014_));
 sky130_fd_sc_hd__a21oi_2 _22340_ (.A1(_07731_),
    .A2(_08013_),
    .B1(_08014_),
    .Y(_08015_));
 sky130_fd_sc_hd__o2bb2ai_2 _22341_ (.A1_N(_08008_),
    .A2_N(_08015_),
    .B1(_08008_),
    .B2(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__a2bb2o_2 _22342_ (.A1_N(_07867_),
    .A2_N(_08016_),
    .B1(_07867_),
    .B2(_08016_),
    .X(_08017_));
 sky130_fd_sc_hd__o22a_2 _22343_ (.A1(_07886_),
    .A2(_07891_),
    .B1(_07885_),
    .B2(_07892_),
    .X(_08018_));
 sky130_fd_sc_hd__o22a_2 _22344_ (.A1(_07912_),
    .A2(_07913_),
    .B1(_07907_),
    .B2(_07914_),
    .X(_08019_));
 sky130_fd_sc_hd__a21oi_2 _22345_ (.A1(_07889_),
    .A2(_07890_),
    .B1(_07888_),
    .Y(_08020_));
 sky130_fd_sc_hd__o21ba_2 _22346_ (.A1(_07903_),
    .A2(_07906_),
    .B1_N(_07905_),
    .X(_08021_));
 sky130_fd_sc_hd__o22a_2 _22347_ (.A1(_07602_),
    .A2(_07009_),
    .B1(_04828_),
    .B2(_07023_),
    .X(_08022_));
 sky130_fd_sc_hd__and4_2 _22348_ (.A(_11620_),
    .B(_11880_),
    .C(_11624_),
    .D(_11877_),
    .X(_08023_));
 sky130_fd_sc_hd__nor2_2 _22349_ (.A(_08022_),
    .B(_08023_),
    .Y(_08024_));
 sky130_fd_sc_hd__nor2_2 _22350_ (.A(_04795_),
    .B(_07160_),
    .Y(_08025_));
 sky130_fd_sc_hd__a2bb2o_2 _22351_ (.A1_N(_08024_),
    .A2_N(_08025_),
    .B1(_08024_),
    .B2(_08025_),
    .X(_08026_));
 sky130_fd_sc_hd__a2bb2o_2 _22352_ (.A1_N(_08021_),
    .A2_N(_08026_),
    .B1(_08021_),
    .B2(_08026_),
    .X(_08027_));
 sky130_fd_sc_hd__a2bb2o_2 _22353_ (.A1_N(_08020_),
    .A2_N(_08027_),
    .B1(_08020_),
    .B2(_08027_),
    .X(_08028_));
 sky130_fd_sc_hd__a2bb2o_2 _22354_ (.A1_N(_08019_),
    .A2_N(_08028_),
    .B1(_08019_),
    .B2(_08028_),
    .X(_08029_));
 sky130_fd_sc_hd__a2bb2o_2 _22355_ (.A1_N(_08018_),
    .A2_N(_08029_),
    .B1(_08018_),
    .B2(_08029_),
    .X(_08030_));
 sky130_fd_sc_hd__o22a_2 _22356_ (.A1(_07884_),
    .A2(_07893_),
    .B1(_07883_),
    .B2(_07894_),
    .X(_08031_));
 sky130_fd_sc_hd__a2bb2o_2 _22357_ (.A1_N(_08030_),
    .A2_N(_08031_),
    .B1(_08030_),
    .B2(_08031_),
    .X(_08032_));
 sky130_fd_sc_hd__a2bb2o_2 _22358_ (.A1_N(_08017_),
    .A2_N(_08032_),
    .B1(_08017_),
    .B2(_08032_),
    .X(_08033_));
 sky130_fd_sc_hd__a2bb2o_2 _22359_ (.A1_N(_08007_),
    .A2_N(_08033_),
    .B1(_08007_),
    .B2(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__a2bb2o_2 _22360_ (.A1_N(_08006_),
    .A2_N(_08034_),
    .B1(_08006_),
    .B2(_08034_),
    .X(_08035_));
 sky130_fd_sc_hd__o22a_2 _22361_ (.A1(_07926_),
    .A2(_07927_),
    .B1(_07915_),
    .B2(_07928_),
    .X(_08036_));
 sky130_fd_sc_hd__o22a_2 _22362_ (.A1(_07933_),
    .A2(_07946_),
    .B1(_07932_),
    .B2(_07947_),
    .X(_08037_));
 sky130_fd_sc_hd__buf_1 _22363_ (.A(_05779_),
    .X(_08038_));
 sky130_fd_sc_hd__o22a_2 _22364_ (.A1(_08038_),
    .A2(_06496_),
    .B1(_04951_),
    .B2(_06624_),
    .X(_08039_));
 sky130_fd_sc_hd__and4_2 _22365_ (.A(_11614_),
    .B(_11888_),
    .C(_11617_),
    .D(_07155_),
    .X(_08040_));
 sky130_fd_sc_hd__nor2_2 _22366_ (.A(_08039_),
    .B(_08040_),
    .Y(_08041_));
 sky130_fd_sc_hd__nor2_2 _22367_ (.A(_04903_),
    .B(_07008_),
    .Y(_08042_));
 sky130_fd_sc_hd__a2bb2o_2 _22368_ (.A1_N(_08041_),
    .A2_N(_08042_),
    .B1(_08041_),
    .B2(_08042_),
    .X(_08043_));
 sky130_fd_sc_hd__or2_2 _22369_ (.A(_07624_),
    .B(_06377_),
    .X(_08044_));
 sky130_fd_sc_hd__o22a_2 _22370_ (.A1(_07626_),
    .A2(_06111_),
    .B1(_05132_),
    .B2(_07173_),
    .X(_08045_));
 sky130_fd_sc_hd__and4_2 _22371_ (.A(_11608_),
    .B(_07038_),
    .C(_11611_),
    .D(_07175_),
    .X(_08046_));
 sky130_fd_sc_hd__or2_2 _22372_ (.A(_08045_),
    .B(_08046_),
    .X(_08047_));
 sky130_fd_sc_hd__a2bb2o_2 _22373_ (.A1_N(_08044_),
    .A2_N(_08047_),
    .B1(_08044_),
    .B2(_08047_),
    .X(_08048_));
 sky130_fd_sc_hd__o21ba_2 _22374_ (.A1(_07908_),
    .A2(_07911_),
    .B1_N(_07910_),
    .X(_08049_));
 sky130_fd_sc_hd__a2bb2o_2 _22375_ (.A1_N(_08048_),
    .A2_N(_08049_),
    .B1(_08048_),
    .B2(_08049_),
    .X(_08050_));
 sky130_fd_sc_hd__a2bb2o_2 _22376_ (.A1_N(_08043_),
    .A2_N(_08050_),
    .B1(_08043_),
    .B2(_08050_),
    .X(_08051_));
 sky130_fd_sc_hd__a21oi_2 _22377_ (.A1(_07921_),
    .A2(_07923_),
    .B1(_07920_),
    .Y(_08052_));
 sky130_fd_sc_hd__o21ba_2 _22378_ (.A1(_07934_),
    .A2(_07937_),
    .B1_N(_07936_),
    .X(_08053_));
 sky130_fd_sc_hd__o22a_2 _22379_ (.A1(_07918_),
    .A2(_05823_),
    .B1(_05389_),
    .B2(_05892_),
    .X(_08054_));
 sky130_fd_sc_hd__and4_2 _22380_ (.A(_11603_),
    .B(_06240_),
    .C(_11606_),
    .D(_11902_),
    .X(_08055_));
 sky130_fd_sc_hd__nor2_2 _22381_ (.A(_08054_),
    .B(_08055_),
    .Y(_08056_));
 sky130_fd_sc_hd__buf_1 _22382_ (.A(_06904_),
    .X(_08057_));
 sky130_fd_sc_hd__nor2_2 _22383_ (.A(_05310_),
    .B(_08057_),
    .Y(_08058_));
 sky130_fd_sc_hd__a2bb2o_2 _22384_ (.A1_N(_08056_),
    .A2_N(_08058_),
    .B1(_08056_),
    .B2(_08058_),
    .X(_08059_));
 sky130_fd_sc_hd__a2bb2o_2 _22385_ (.A1_N(_08053_),
    .A2_N(_08059_),
    .B1(_08053_),
    .B2(_08059_),
    .X(_08060_));
 sky130_fd_sc_hd__a2bb2o_2 _22386_ (.A1_N(_08052_),
    .A2_N(_08060_),
    .B1(_08052_),
    .B2(_08060_),
    .X(_08061_));
 sky130_fd_sc_hd__o22a_2 _22387_ (.A1(_07917_),
    .A2(_07924_),
    .B1(_07916_),
    .B2(_07925_),
    .X(_08062_));
 sky130_fd_sc_hd__a2bb2o_2 _22388_ (.A1_N(_08061_),
    .A2_N(_08062_),
    .B1(_08061_),
    .B2(_08062_),
    .X(_08063_));
 sky130_fd_sc_hd__a2bb2o_2 _22389_ (.A1_N(_08051_),
    .A2_N(_08063_),
    .B1(_08051_),
    .B2(_08063_),
    .X(_08064_));
 sky130_fd_sc_hd__a2bb2o_2 _22390_ (.A1_N(_08037_),
    .A2_N(_08064_),
    .B1(_08037_),
    .B2(_08064_),
    .X(_08065_));
 sky130_fd_sc_hd__a2bb2o_2 _22391_ (.A1_N(_08036_),
    .A2_N(_08065_),
    .B1(_08036_),
    .B2(_08065_),
    .X(_08066_));
 sky130_fd_sc_hd__o22a_2 _22392_ (.A1(_07943_),
    .A2(_07944_),
    .B1(_07938_),
    .B2(_07945_),
    .X(_08067_));
 sky130_fd_sc_hd__o22a_2 _22393_ (.A1(_07950_),
    .A2(_07955_),
    .B1(_07949_),
    .B2(_07956_),
    .X(_08068_));
 sky130_fd_sc_hd__or2_2 _22394_ (.A(_05562_),
    .B(_05716_),
    .X(_08069_));
 sky130_fd_sc_hd__o22a_2 _22395_ (.A1(_07359_),
    .A2(_06257_),
    .B1(_05659_),
    .B2(_06254_),
    .X(_08070_));
 sky130_fd_sc_hd__and4_2 _22396_ (.A(_11593_),
    .B(_06392_),
    .C(_11598_),
    .D(_06393_),
    .X(_08071_));
 sky130_fd_sc_hd__or2_2 _22397_ (.A(_08070_),
    .B(_08071_),
    .X(_08072_));
 sky130_fd_sc_hd__a2bb2o_2 _22398_ (.A1_N(_08069_),
    .A2_N(_08072_),
    .B1(_08069_),
    .B2(_08072_),
    .X(_08073_));
 sky130_fd_sc_hd__or2_2 _22399_ (.A(_07656_),
    .B(_05828_),
    .X(_08074_));
 sky130_fd_sc_hd__o22a_2 _22400_ (.A1(_07658_),
    .A2(_05334_),
    .B1(_06034_),
    .B2(_05420_),
    .X(_08075_));
 sky130_fd_sc_hd__and4_2 _22401_ (.A(_07515_),
    .B(_07509_),
    .C(_07516_),
    .D(_06016_),
    .X(_08076_));
 sky130_fd_sc_hd__or2_2 _22402_ (.A(_08075_),
    .B(_08076_),
    .X(_08077_));
 sky130_fd_sc_hd__a2bb2o_2 _22403_ (.A1_N(_08074_),
    .A2_N(_08077_),
    .B1(_08074_),
    .B2(_08077_),
    .X(_08078_));
 sky130_fd_sc_hd__o21ba_2 _22404_ (.A1(_07939_),
    .A2(_07942_),
    .B1_N(_07941_),
    .X(_08079_));
 sky130_fd_sc_hd__a2bb2o_2 _22405_ (.A1_N(_08078_),
    .A2_N(_08079_),
    .B1(_08078_),
    .B2(_08079_),
    .X(_08080_));
 sky130_fd_sc_hd__a2bb2o_2 _22406_ (.A1_N(_08073_),
    .A2_N(_08080_),
    .B1(_08073_),
    .B2(_08080_),
    .X(_08081_));
 sky130_fd_sc_hd__a2bb2o_2 _22407_ (.A1_N(_08068_),
    .A2_N(_08081_),
    .B1(_08068_),
    .B2(_08081_),
    .X(_08082_));
 sky130_fd_sc_hd__a2bb2o_2 _22408_ (.A1_N(_08067_),
    .A2_N(_08082_),
    .B1(_08067_),
    .B2(_08082_),
    .X(_08083_));
 sky130_fd_sc_hd__o21ba_2 _22409_ (.A1(_07951_),
    .A2(_07954_),
    .B1_N(_07953_),
    .X(_08084_));
 sky130_fd_sc_hd__o21ba_2 _22410_ (.A1(_07958_),
    .A2(_07961_),
    .B1_N(_07960_),
    .X(_08085_));
 sky130_fd_sc_hd__or2_2 _22411_ (.A(_07376_),
    .B(_05247_),
    .X(_08086_));
 sky130_fd_sc_hd__o22a_2 _22412_ (.A1(_07378_),
    .A2(_05530_),
    .B1(_07379_),
    .B2(_05740_),
    .X(_08087_));
 sky130_fd_sc_hd__and4_2 _22413_ (.A(_07240_),
    .B(_11927_),
    .C(_07672_),
    .D(_05745_),
    .X(_08088_));
 sky130_fd_sc_hd__or2_2 _22414_ (.A(_08087_),
    .B(_08088_),
    .X(_08089_));
 sky130_fd_sc_hd__a2bb2o_2 _22415_ (.A1_N(_08086_),
    .A2_N(_08089_),
    .B1(_08086_),
    .B2(_08089_),
    .X(_08090_));
 sky130_fd_sc_hd__a2bb2o_2 _22416_ (.A1_N(_08085_),
    .A2_N(_08090_),
    .B1(_08085_),
    .B2(_08090_),
    .X(_08091_));
 sky130_fd_sc_hd__a2bb2o_2 _22417_ (.A1_N(_08084_),
    .A2_N(_08091_),
    .B1(_08084_),
    .B2(_08091_),
    .X(_08092_));
 sky130_fd_sc_hd__or2_2 _22418_ (.A(_06686_),
    .B(_05164_),
    .X(_08093_));
 sky130_fd_sc_hd__o22a_2 _22419_ (.A1(_07387_),
    .A2(_05273_),
    .B1(_06829_),
    .B2(_05943_),
    .X(_08094_));
 sky130_fd_sc_hd__and4_2 _22420_ (.A(_07538_),
    .B(_11934_),
    .C(_07539_),
    .D(_05781_),
    .X(_08095_));
 sky130_fd_sc_hd__or2_2 _22421_ (.A(_08094_),
    .B(_08095_),
    .X(_08096_));
 sky130_fd_sc_hd__a2bb2o_2 _22422_ (.A1_N(_08093_),
    .A2_N(_08096_),
    .B1(_08093_),
    .B2(_08096_),
    .X(_08097_));
 sky130_fd_sc_hd__buf_1 _22423_ (.A(_07099_),
    .X(_08098_));
 sky130_fd_sc_hd__or2_2 _22424_ (.A(_08098_),
    .B(_05191_),
    .X(_08099_));
 sky130_fd_sc_hd__buf_1 _22425_ (.A(\pcpi_mul.rs2[31] ),
    .X(_08100_));
 sky130_fd_sc_hd__and4_2 _22426_ (.A(_07830_),
    .B(_05194_),
    .C(_08100_),
    .D(_05198_),
    .X(_08101_));
 sky130_fd_sc_hd__o22a_2 _22427_ (.A1(_07832_),
    .A2(_05197_),
    .B1(_07965_),
    .B2(_05195_),
    .X(_08102_));
 sky130_fd_sc_hd__or2_2 _22428_ (.A(_08101_),
    .B(_08102_),
    .X(_08103_));
 sky130_fd_sc_hd__a2bb2o_2 _22429_ (.A1_N(_08099_),
    .A2_N(_08103_),
    .B1(_08099_),
    .B2(_08103_),
    .X(_08104_));
 sky130_fd_sc_hd__o21ba_2 _22430_ (.A1(_07963_),
    .A2(_07967_),
    .B1_N(_07964_),
    .X(_08105_));
 sky130_fd_sc_hd__a2bb2o_2 _22431_ (.A1_N(_08104_),
    .A2_N(_08105_),
    .B1(_08104_),
    .B2(_08105_),
    .X(_08106_));
 sky130_fd_sc_hd__a2bb2o_2 _22432_ (.A1_N(_08097_),
    .A2_N(_08106_),
    .B1(_08097_),
    .B2(_08106_),
    .X(_08107_));
 sky130_fd_sc_hd__o22a_2 _22433_ (.A1(_07968_),
    .A2(_07969_),
    .B1(_07962_),
    .B2(_07970_),
    .X(_08108_));
 sky130_fd_sc_hd__a2bb2o_2 _22434_ (.A1_N(_08107_),
    .A2_N(_08108_),
    .B1(_08107_),
    .B2(_08108_),
    .X(_08109_));
 sky130_fd_sc_hd__a2bb2o_2 _22435_ (.A1_N(_08092_),
    .A2_N(_08109_),
    .B1(_08092_),
    .B2(_08109_),
    .X(_08110_));
 sky130_fd_sc_hd__o22a_2 _22436_ (.A1(_07971_),
    .A2(_07972_),
    .B1(_07957_),
    .B2(_07973_),
    .X(_08111_));
 sky130_fd_sc_hd__a2bb2o_2 _22437_ (.A1_N(_08110_),
    .A2_N(_08111_),
    .B1(_08110_),
    .B2(_08111_),
    .X(_08112_));
 sky130_fd_sc_hd__a2bb2o_2 _22438_ (.A1_N(_08083_),
    .A2_N(_08112_),
    .B1(_08083_),
    .B2(_08112_),
    .X(_08113_));
 sky130_fd_sc_hd__o22a_2 _22439_ (.A1(_07974_),
    .A2(_07975_),
    .B1(_07948_),
    .B2(_07976_),
    .X(_08114_));
 sky130_fd_sc_hd__a2bb2o_2 _22440_ (.A1_N(_08113_),
    .A2_N(_08114_),
    .B1(_08113_),
    .B2(_08114_),
    .X(_08115_));
 sky130_fd_sc_hd__a2bb2o_2 _22441_ (.A1_N(_08066_),
    .A2_N(_08115_),
    .B1(_08066_),
    .B2(_08115_),
    .X(_08116_));
 sky130_fd_sc_hd__o22a_2 _22442_ (.A1(_07977_),
    .A2(_07978_),
    .B1(_07931_),
    .B2(_07979_),
    .X(_08117_));
 sky130_fd_sc_hd__a2bb2o_2 _22443_ (.A1_N(_08116_),
    .A2_N(_08117_),
    .B1(_08116_),
    .B2(_08117_),
    .X(_08118_));
 sky130_fd_sc_hd__a2bb2o_2 _22444_ (.A1_N(_08035_),
    .A2_N(_08118_),
    .B1(_08035_),
    .B2(_08118_),
    .X(_08119_));
 sky130_fd_sc_hd__o22a_2 _22445_ (.A1(_07980_),
    .A2(_07981_),
    .B1(_07900_),
    .B2(_07982_),
    .X(_08120_));
 sky130_fd_sc_hd__a2bb2o_2 _22446_ (.A1_N(_08119_),
    .A2_N(_08120_),
    .B1(_08119_),
    .B2(_08120_),
    .X(_08121_));
 sky130_fd_sc_hd__a2bb2o_2 _22447_ (.A1_N(_08005_),
    .A2_N(_08121_),
    .B1(_08005_),
    .B2(_08121_),
    .X(_08122_));
 sky130_fd_sc_hd__o22a_2 _22448_ (.A1(_07983_),
    .A2(_07984_),
    .B1(_07863_),
    .B2(_07985_),
    .X(_08123_));
 sky130_fd_sc_hd__a2bb2o_2 _22449_ (.A1_N(_08122_),
    .A2_N(_08123_),
    .B1(_08122_),
    .B2(_08123_),
    .X(_08124_));
 sky130_fd_sc_hd__a2bb2o_2 _22450_ (.A1_N(_07862_),
    .A2_N(_08124_),
    .B1(_07862_),
    .B2(_08124_),
    .X(_08125_));
 sky130_fd_sc_hd__or2_2 _22451_ (.A(_08000_),
    .B(_08125_),
    .X(_08126_));
 sky130_fd_sc_hd__a21bo_2 _22452_ (.A1(_08000_),
    .A2(_08125_),
    .B1_N(_08126_),
    .X(_08127_));
 sky130_fd_sc_hd__o21ai_2 _22453_ (.A1(_07992_),
    .A2(_07998_),
    .B1(_07991_),
    .Y(_08128_));
 sky130_fd_sc_hd__a2bb2o_2 _22454_ (.A1_N(_08127_),
    .A2_N(_08128_),
    .B1(_08127_),
    .B2(_08128_),
    .X(_02656_));
 sky130_fd_sc_hd__o22a_2 _22455_ (.A1(_08007_),
    .A2(_08033_),
    .B1(_08006_),
    .B2(_08034_),
    .X(_08129_));
 sky130_fd_sc_hd__o22a_2 _22456_ (.A1(_08008_),
    .A2(_08015_),
    .B1(_08002_),
    .B2(_08016_),
    .X(_08130_));
 sky130_fd_sc_hd__or2_2 _22457_ (.A(_08129_),
    .B(_08130_),
    .X(_08131_));
 sky130_fd_sc_hd__a21bo_2 _22458_ (.A1(_08129_),
    .A2(_08130_),
    .B1_N(_08131_),
    .X(_08132_));
 sky130_fd_sc_hd__o22a_2 _22459_ (.A1(_08030_),
    .A2(_08031_),
    .B1(_08017_),
    .B2(_08032_),
    .X(_08133_));
 sky130_fd_sc_hd__o22a_2 _22460_ (.A1(_08037_),
    .A2(_08064_),
    .B1(_08036_),
    .B2(_08065_),
    .X(_08134_));
 sky130_fd_sc_hd__or2_2 _22461_ (.A(_07447_),
    .B(_08010_),
    .X(_08135_));
 sky130_vsdinv _22462_ (.A(_08135_),
    .Y(_08136_));
 sky130_fd_sc_hd__o32a_2 _22463_ (.A1(_07731_),
    .A2(_08013_),
    .A3(_08135_),
    .B1(_08014_),
    .B2(_08136_),
    .X(_08137_));
 sky130_fd_sc_hd__a2bb2o_2 _22464_ (.A1_N(_08002_),
    .A2_N(_08137_),
    .B1(_08002_),
    .B2(_08137_),
    .X(_08138_));
 sky130_fd_sc_hd__o22a_2 _22465_ (.A1(_08021_),
    .A2(_08026_),
    .B1(_08020_),
    .B2(_08027_),
    .X(_08139_));
 sky130_fd_sc_hd__o22a_2 _22466_ (.A1(_08048_),
    .A2(_08049_),
    .B1(_08043_),
    .B2(_08050_),
    .X(_08140_));
 sky130_fd_sc_hd__a21oi_2 _22467_ (.A1(_08024_),
    .A2(_08025_),
    .B1(_08023_),
    .Y(_08141_));
 sky130_fd_sc_hd__a21oi_2 _22468_ (.A1(_08041_),
    .A2(_08042_),
    .B1(_08040_),
    .Y(_08142_));
 sky130_fd_sc_hd__o22a_2 _22469_ (.A1(_05193_),
    .A2(_07022_),
    .B1(_04827_),
    .B2(_07732_),
    .X(_08143_));
 sky130_fd_sc_hd__and4_2 _22470_ (.A(_11619_),
    .B(_11876_),
    .C(_11623_),
    .D(\pcpi_mul.rs1[31] ),
    .X(_08144_));
 sky130_fd_sc_hd__or2_2 _22471_ (.A(_08143_),
    .B(_08144_),
    .X(_08145_));
 sky130_vsdinv _22472_ (.A(_08145_),
    .Y(_08146_));
 sky130_fd_sc_hd__or2_2 _22473_ (.A(_10585_),
    .B(_04793_),
    .X(_08147_));
 sky130_fd_sc_hd__buf_1 _22474_ (.A(_08147_),
    .X(_08148_));
 sky130_fd_sc_hd__a32o_2 _22475_ (.A1(_07869_),
    .A2(\pcpi_mul.rs2[6] ),
    .A3(_08146_),
    .B1(_08145_),
    .B2(_08148_),
    .X(_08149_));
 sky130_fd_sc_hd__a2bb2o_2 _22476_ (.A1_N(_08142_),
    .A2_N(_08149_),
    .B1(_08142_),
    .B2(_08149_),
    .X(_08150_));
 sky130_fd_sc_hd__a2bb2o_2 _22477_ (.A1_N(_08141_),
    .A2_N(_08150_),
    .B1(_08141_),
    .B2(_08150_),
    .X(_08151_));
 sky130_fd_sc_hd__a2bb2o_2 _22478_ (.A1_N(_08140_),
    .A2_N(_08151_),
    .B1(_08140_),
    .B2(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__a2bb2o_2 _22479_ (.A1_N(_08139_),
    .A2_N(_08152_),
    .B1(_08139_),
    .B2(_08152_),
    .X(_08153_));
 sky130_fd_sc_hd__o22a_2 _22480_ (.A1(_08019_),
    .A2(_08028_),
    .B1(_08018_),
    .B2(_08029_),
    .X(_08154_));
 sky130_fd_sc_hd__a2bb2o_2 _22481_ (.A1_N(_08153_),
    .A2_N(_08154_),
    .B1(_08153_),
    .B2(_08154_),
    .X(_08155_));
 sky130_fd_sc_hd__a2bb2o_2 _22482_ (.A1_N(_08138_),
    .A2_N(_08155_),
    .B1(_08138_),
    .B2(_08155_),
    .X(_08156_));
 sky130_fd_sc_hd__a2bb2o_2 _22483_ (.A1_N(_08134_),
    .A2_N(_08156_),
    .B1(_08134_),
    .B2(_08156_),
    .X(_08157_));
 sky130_fd_sc_hd__a2bb2o_2 _22484_ (.A1_N(_08133_),
    .A2_N(_08157_),
    .B1(_08133_),
    .B2(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__o22a_2 _22485_ (.A1(_08061_),
    .A2(_08062_),
    .B1(_08051_),
    .B2(_08063_),
    .X(_08159_));
 sky130_fd_sc_hd__o22a_2 _22486_ (.A1(_08068_),
    .A2(_08081_),
    .B1(_08067_),
    .B2(_08082_),
    .X(_08160_));
 sky130_fd_sc_hd__o22a_2 _22487_ (.A1(_08038_),
    .A2(_06624_),
    .B1(_04951_),
    .B2(_07007_),
    .X(_08161_));
 sky130_fd_sc_hd__and4_2 _22488_ (.A(_11614_),
    .B(_07155_),
    .C(_11617_),
    .D(_11882_),
    .X(_08162_));
 sky130_fd_sc_hd__nor2_2 _22489_ (.A(_08161_),
    .B(_08162_),
    .Y(_08163_));
 sky130_fd_sc_hd__nor2_2 _22490_ (.A(_04903_),
    .B(_07010_),
    .Y(_08164_));
 sky130_fd_sc_hd__a2bb2o_2 _22491_ (.A1_N(_08163_),
    .A2_N(_08164_),
    .B1(_08163_),
    .B2(_08164_),
    .X(_08165_));
 sky130_fd_sc_hd__or2_2 _22492_ (.A(_07624_),
    .B(_06743_),
    .X(_08166_));
 sky130_fd_sc_hd__o22a_2 _22493_ (.A1(_07626_),
    .A2(_07173_),
    .B1(_07481_),
    .B2(_06376_),
    .X(_08167_));
 sky130_fd_sc_hd__and4_2 _22494_ (.A(_11608_),
    .B(_07175_),
    .C(_11611_),
    .D(_11892_),
    .X(_08168_));
 sky130_fd_sc_hd__or2_2 _22495_ (.A(_08167_),
    .B(_08168_),
    .X(_08169_));
 sky130_fd_sc_hd__a2bb2o_2 _22496_ (.A1_N(_08166_),
    .A2_N(_08169_),
    .B1(_08166_),
    .B2(_08169_),
    .X(_08170_));
 sky130_fd_sc_hd__o21ba_2 _22497_ (.A1(_08044_),
    .A2(_08047_),
    .B1_N(_08046_),
    .X(_08171_));
 sky130_fd_sc_hd__a2bb2o_2 _22498_ (.A1_N(_08170_),
    .A2_N(_08171_),
    .B1(_08170_),
    .B2(_08171_),
    .X(_08172_));
 sky130_fd_sc_hd__a2bb2o_2 _22499_ (.A1_N(_08165_),
    .A2_N(_08172_),
    .B1(_08165_),
    .B2(_08172_),
    .X(_08173_));
 sky130_fd_sc_hd__a21oi_2 _22500_ (.A1(_08056_),
    .A2(_08058_),
    .B1(_08055_),
    .Y(_08174_));
 sky130_fd_sc_hd__o21ba_2 _22501_ (.A1(_08069_),
    .A2(_08072_),
    .B1_N(_08071_),
    .X(_08175_));
 sky130_fd_sc_hd__buf_1 _22502_ (.A(_05388_),
    .X(_08176_));
 sky130_fd_sc_hd__o22a_2 _22503_ (.A1(_07918_),
    .A2(_06501_),
    .B1(_08176_),
    .B2(_06904_),
    .X(_08177_));
 sky130_fd_sc_hd__and4_2 _22504_ (.A(_11603_),
    .B(_11902_),
    .C(_11606_),
    .D(_06499_),
    .X(_08178_));
 sky130_fd_sc_hd__nor2_2 _22505_ (.A(_08177_),
    .B(_08178_),
    .Y(_08179_));
 sky130_fd_sc_hd__nor2_2 _22506_ (.A(_07922_),
    .B(_06112_),
    .Y(_08180_));
 sky130_fd_sc_hd__a2bb2o_2 _22507_ (.A1_N(_08179_),
    .A2_N(_08180_),
    .B1(_08179_),
    .B2(_08180_),
    .X(_08181_));
 sky130_fd_sc_hd__a2bb2o_2 _22508_ (.A1_N(_08175_),
    .A2_N(_08181_),
    .B1(_08175_),
    .B2(_08181_),
    .X(_08182_));
 sky130_fd_sc_hd__a2bb2o_2 _22509_ (.A1_N(_08174_),
    .A2_N(_08182_),
    .B1(_08174_),
    .B2(_08182_),
    .X(_08183_));
 sky130_fd_sc_hd__o22a_2 _22510_ (.A1(_08053_),
    .A2(_08059_),
    .B1(_08052_),
    .B2(_08060_),
    .X(_08184_));
 sky130_fd_sc_hd__a2bb2o_2 _22511_ (.A1_N(_08183_),
    .A2_N(_08184_),
    .B1(_08183_),
    .B2(_08184_),
    .X(_08185_));
 sky130_fd_sc_hd__a2bb2o_2 _22512_ (.A1_N(_08173_),
    .A2_N(_08185_),
    .B1(_08173_),
    .B2(_08185_),
    .X(_08186_));
 sky130_fd_sc_hd__a2bb2o_2 _22513_ (.A1_N(_08160_),
    .A2_N(_08186_),
    .B1(_08160_),
    .B2(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__a2bb2o_2 _22514_ (.A1_N(_08159_),
    .A2_N(_08187_),
    .B1(_08159_),
    .B2(_08187_),
    .X(_08188_));
 sky130_fd_sc_hd__o22a_2 _22515_ (.A1(_08078_),
    .A2(_08079_),
    .B1(_08073_),
    .B2(_08080_),
    .X(_08189_));
 sky130_fd_sc_hd__o22a_2 _22516_ (.A1(_08085_),
    .A2(_08090_),
    .B1(_08084_),
    .B2(_08091_),
    .X(_08190_));
 sky130_fd_sc_hd__or2_2 _22517_ (.A(_06700_),
    .B(_06237_),
    .X(_08191_));
 sky130_fd_sc_hd__o22a_2 _22518_ (.A1(_07359_),
    .A2(_06254_),
    .B1(_05662_),
    .B2(_05715_),
    .X(_08192_));
 sky130_fd_sc_hd__and4_2 _22519_ (.A(_06703_),
    .B(_06393_),
    .C(_11598_),
    .D(_11908_),
    .X(_08193_));
 sky130_fd_sc_hd__or2_2 _22520_ (.A(_08192_),
    .B(_08193_),
    .X(_08194_));
 sky130_fd_sc_hd__a2bb2o_2 _22521_ (.A1_N(_08191_),
    .A2_N(_08194_),
    .B1(_08191_),
    .B2(_08194_),
    .X(_08195_));
 sky130_fd_sc_hd__or2_2 _22522_ (.A(_07656_),
    .B(_05510_),
    .X(_08196_));
 sky130_fd_sc_hd__o22a_2 _22523_ (.A1(_07658_),
    .A2(_06014_),
    .B1(_06030_),
    .B2(_06134_),
    .X(_08197_));
 sky130_fd_sc_hd__and4_2 _22524_ (.A(_07515_),
    .B(_06016_),
    .C(_07516_),
    .D(_06138_),
    .X(_08198_));
 sky130_fd_sc_hd__or2_2 _22525_ (.A(_08197_),
    .B(_08198_),
    .X(_08199_));
 sky130_fd_sc_hd__a2bb2o_2 _22526_ (.A1_N(_08196_),
    .A2_N(_08199_),
    .B1(_08196_),
    .B2(_08199_),
    .X(_08200_));
 sky130_fd_sc_hd__o21ba_2 _22527_ (.A1(_08074_),
    .A2(_08077_),
    .B1_N(_08076_),
    .X(_08201_));
 sky130_fd_sc_hd__a2bb2o_2 _22528_ (.A1_N(_08200_),
    .A2_N(_08201_),
    .B1(_08200_),
    .B2(_08201_),
    .X(_08202_));
 sky130_fd_sc_hd__a2bb2o_2 _22529_ (.A1_N(_08195_),
    .A2_N(_08202_),
    .B1(_08195_),
    .B2(_08202_),
    .X(_08203_));
 sky130_fd_sc_hd__a2bb2o_2 _22530_ (.A1_N(_08190_),
    .A2_N(_08203_),
    .B1(_08190_),
    .B2(_08203_),
    .X(_08204_));
 sky130_fd_sc_hd__a2bb2o_2 _22531_ (.A1_N(_08189_),
    .A2_N(_08204_),
    .B1(_08189_),
    .B2(_08204_),
    .X(_08205_));
 sky130_fd_sc_hd__o21ba_2 _22532_ (.A1(_08086_),
    .A2(_08089_),
    .B1_N(_08088_),
    .X(_08206_));
 sky130_fd_sc_hd__o21ba_2 _22533_ (.A1(_08093_),
    .A2(_08096_),
    .B1_N(_08095_),
    .X(_08207_));
 sky130_fd_sc_hd__or2_2 _22534_ (.A(_07376_),
    .B(_05335_),
    .X(_08208_));
 sky130_fd_sc_hd__o22a_2 _22535_ (.A1(_07378_),
    .A2(_05157_),
    .B1(_07379_),
    .B2(_05246_),
    .X(_08209_));
 sky130_fd_sc_hd__and4_2 _22536_ (.A(_07240_),
    .B(_05745_),
    .C(_11580_),
    .D(_05848_),
    .X(_08210_));
 sky130_fd_sc_hd__or2_2 _22537_ (.A(_08209_),
    .B(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__a2bb2o_2 _22538_ (.A1_N(_08208_),
    .A2_N(_08211_),
    .B1(_08208_),
    .B2(_08211_),
    .X(_08212_));
 sky130_fd_sc_hd__a2bb2o_2 _22539_ (.A1_N(_08207_),
    .A2_N(_08212_),
    .B1(_08207_),
    .B2(_08212_),
    .X(_08213_));
 sky130_fd_sc_hd__a2bb2o_2 _22540_ (.A1_N(_08206_),
    .A2_N(_08213_),
    .B1(_08206_),
    .B2(_08213_),
    .X(_08214_));
 sky130_fd_sc_hd__or2_2 _22541_ (.A(_06685_),
    .B(_05155_),
    .X(_08215_));
 sky130_fd_sc_hd__o22a_2 _22542_ (.A1(_07387_),
    .A2(_06429_),
    .B1(_06829_),
    .B2(_06180_),
    .X(_08216_));
 sky130_fd_sc_hd__and4_2 _22543_ (.A(_11566_),
    .B(_05781_),
    .C(_07539_),
    .D(_06184_),
    .X(_08217_));
 sky130_fd_sc_hd__or2_2 _22544_ (.A(_08216_),
    .B(_08217_),
    .X(_08218_));
 sky130_fd_sc_hd__a2bb2o_2 _22545_ (.A1_N(_08215_),
    .A2_N(_08218_),
    .B1(_08215_),
    .B2(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__or2_2 _22546_ (.A(_07828_),
    .B(_06568_),
    .X(_08220_));
 sky130_fd_sc_hd__and4_2 _22547_ (.A(_07830_),
    .B(_05398_),
    .C(_11560_),
    .D(_05280_),
    .X(_08221_));
 sky130_fd_sc_hd__o22a_2 _22548_ (.A1(_07832_),
    .A2(_05198_),
    .B1(_07247_),
    .B2(_05190_),
    .X(_08222_));
 sky130_fd_sc_hd__or2_2 _22549_ (.A(_08221_),
    .B(_08222_),
    .X(_08223_));
 sky130_fd_sc_hd__a2bb2o_2 _22550_ (.A1_N(_08220_),
    .A2_N(_08223_),
    .B1(_08220_),
    .B2(_08223_),
    .X(_08224_));
 sky130_fd_sc_hd__o21ba_2 _22551_ (.A1(_08099_),
    .A2(_08103_),
    .B1_N(_08101_),
    .X(_08225_));
 sky130_fd_sc_hd__a2bb2o_2 _22552_ (.A1_N(_08224_),
    .A2_N(_08225_),
    .B1(_08224_),
    .B2(_08225_),
    .X(_08226_));
 sky130_fd_sc_hd__a2bb2o_2 _22553_ (.A1_N(_08219_),
    .A2_N(_08226_),
    .B1(_08219_),
    .B2(_08226_),
    .X(_08227_));
 sky130_fd_sc_hd__o22a_2 _22554_ (.A1(_08104_),
    .A2(_08105_),
    .B1(_08097_),
    .B2(_08106_),
    .X(_08228_));
 sky130_fd_sc_hd__a2bb2o_2 _22555_ (.A1_N(_08227_),
    .A2_N(_08228_),
    .B1(_08227_),
    .B2(_08228_),
    .X(_08229_));
 sky130_fd_sc_hd__a2bb2o_2 _22556_ (.A1_N(_08214_),
    .A2_N(_08229_),
    .B1(_08214_),
    .B2(_08229_),
    .X(_08230_));
 sky130_fd_sc_hd__o22a_2 _22557_ (.A1(_08107_),
    .A2(_08108_),
    .B1(_08092_),
    .B2(_08109_),
    .X(_08231_));
 sky130_fd_sc_hd__a2bb2o_2 _22558_ (.A1_N(_08230_),
    .A2_N(_08231_),
    .B1(_08230_),
    .B2(_08231_),
    .X(_08232_));
 sky130_fd_sc_hd__a2bb2o_2 _22559_ (.A1_N(_08205_),
    .A2_N(_08232_),
    .B1(_08205_),
    .B2(_08232_),
    .X(_08233_));
 sky130_fd_sc_hd__o22a_2 _22560_ (.A1(_08110_),
    .A2(_08111_),
    .B1(_08083_),
    .B2(_08112_),
    .X(_08234_));
 sky130_fd_sc_hd__a2bb2o_2 _22561_ (.A1_N(_08233_),
    .A2_N(_08234_),
    .B1(_08233_),
    .B2(_08234_),
    .X(_08235_));
 sky130_fd_sc_hd__a2bb2o_2 _22562_ (.A1_N(_08188_),
    .A2_N(_08235_),
    .B1(_08188_),
    .B2(_08235_),
    .X(_08236_));
 sky130_fd_sc_hd__o22a_2 _22563_ (.A1(_08113_),
    .A2(_08114_),
    .B1(_08066_),
    .B2(_08115_),
    .X(_08237_));
 sky130_fd_sc_hd__a2bb2o_2 _22564_ (.A1_N(_08236_),
    .A2_N(_08237_),
    .B1(_08236_),
    .B2(_08237_),
    .X(_08238_));
 sky130_fd_sc_hd__a2bb2o_2 _22565_ (.A1_N(_08158_),
    .A2_N(_08238_),
    .B1(_08158_),
    .B2(_08238_),
    .X(_08239_));
 sky130_fd_sc_hd__o22a_2 _22566_ (.A1(_08116_),
    .A2(_08117_),
    .B1(_08035_),
    .B2(_08118_),
    .X(_08240_));
 sky130_fd_sc_hd__a2bb2o_2 _22567_ (.A1_N(_08239_),
    .A2_N(_08240_),
    .B1(_08239_),
    .B2(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__a2bb2o_2 _22568_ (.A1_N(_08132_),
    .A2_N(_08241_),
    .B1(_08132_),
    .B2(_08241_),
    .X(_08242_));
 sky130_fd_sc_hd__o22a_2 _22569_ (.A1(_08119_),
    .A2(_08120_),
    .B1(_08005_),
    .B2(_08121_),
    .X(_08243_));
 sky130_fd_sc_hd__a2bb2o_2 _22570_ (.A1_N(_08242_),
    .A2_N(_08243_),
    .B1(_08242_),
    .B2(_08243_),
    .X(_08244_));
 sky130_fd_sc_hd__a2bb2o_2 _22571_ (.A1_N(_08004_),
    .A2_N(_08244_),
    .B1(_08004_),
    .B2(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__o22a_2 _22572_ (.A1(_08122_),
    .A2(_08123_),
    .B1(_07862_),
    .B2(_08124_),
    .X(_08246_));
 sky130_fd_sc_hd__or2_2 _22573_ (.A(_08245_),
    .B(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__a21bo_2 _22574_ (.A1(_08245_),
    .A2(_08246_),
    .B1_N(_08247_),
    .X(_08248_));
 sky130_fd_sc_hd__a22o_2 _22575_ (.A1(_08000_),
    .A2(_08125_),
    .B1(_07991_),
    .B2(_08126_),
    .X(_08249_));
 sky130_fd_sc_hd__o31a_2 _22576_ (.A1(_07992_),
    .A2(_08127_),
    .A3(_07998_),
    .B1(_08249_),
    .X(_08250_));
 sky130_fd_sc_hd__a2bb2oi_2 _22577_ (.A1_N(_08248_),
    .A2_N(_08250_),
    .B1(_08248_),
    .B2(_08250_),
    .Y(_02657_));
 sky130_fd_sc_hd__o22a_2 _22578_ (.A1(_08242_),
    .A2(_08243_),
    .B1(_08004_),
    .B2(_08244_),
    .X(_08251_));
 sky130_fd_sc_hd__o22a_2 _22579_ (.A1(_08134_),
    .A2(_08156_),
    .B1(_08133_),
    .B2(_08157_),
    .X(_08252_));
 sky130_fd_sc_hd__or3_2 _22580_ (.A(_04539_),
    .B(_08009_),
    .C(_07730_),
    .X(_08253_));
 sky130_fd_sc_hd__o21a_2 _22581_ (.A1(_08002_),
    .A2(_08137_),
    .B1(_08253_),
    .X(_08254_));
 sky130_fd_sc_hd__or2_2 _22582_ (.A(_08252_),
    .B(_08254_),
    .X(_08255_));
 sky130_fd_sc_hd__a21bo_2 _22583_ (.A1(_08252_),
    .A2(_08254_),
    .B1_N(_08255_),
    .X(_08256_));
 sky130_fd_sc_hd__o22a_2 _22584_ (.A1(_08153_),
    .A2(_08154_),
    .B1(_08138_),
    .B2(_08155_),
    .X(_08257_));
 sky130_fd_sc_hd__o22a_2 _22585_ (.A1(_08160_),
    .A2(_08186_),
    .B1(_08159_),
    .B2(_08187_),
    .X(_08258_));
 sky130_fd_sc_hd__a21bo_2 _22586_ (.A1(_07730_),
    .A2(_08136_),
    .B1_N(_08253_),
    .X(_08259_));
 sky130_fd_sc_hd__a2bb2o_2 _22587_ (.A1_N(_07867_),
    .A2_N(_08259_),
    .B1(_07866_),
    .B2(_08259_),
    .X(_08260_));
 sky130_fd_sc_hd__buf_1 _22588_ (.A(_08260_),
    .X(_08261_));
 sky130_fd_sc_hd__o22a_2 _22589_ (.A1(_08142_),
    .A2(_08149_),
    .B1(_08141_),
    .B2(_08150_),
    .X(_08262_));
 sky130_fd_sc_hd__o22a_2 _22590_ (.A1(_08170_),
    .A2(_08171_),
    .B1(_08165_),
    .B2(_08172_),
    .X(_08263_));
 sky130_fd_sc_hd__o21ba_2 _22591_ (.A1(_08145_),
    .A2(_08148_),
    .B1_N(_08144_),
    .X(_08264_));
 sky130_fd_sc_hd__a21oi_2 _22592_ (.A1(_08163_),
    .A2(_08164_),
    .B1(_08162_),
    .Y(_08265_));
 sky130_fd_sc_hd__buf_1 _22593_ (.A(_07732_),
    .X(_08266_));
 sky130_fd_sc_hd__nor2_2 _22594_ (.A(_07602_),
    .B(_08266_),
    .Y(_08267_));
 sky130_fd_sc_hd__or2_2 _22595_ (.A(_10584_),
    .B(_04825_),
    .X(_08268_));
 sky130_vsdinv _22596_ (.A(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__a2bb2o_2 _22597_ (.A1_N(_08267_),
    .A2_N(_08269_),
    .B1(_08267_),
    .B2(_08269_),
    .X(_08270_));
 sky130_fd_sc_hd__a2bb2o_2 _22598_ (.A1_N(_08148_),
    .A2_N(_08270_),
    .B1(_08148_),
    .B2(_08270_),
    .X(_08271_));
 sky130_fd_sc_hd__a2bb2o_2 _22599_ (.A1_N(_08265_),
    .A2_N(_08271_),
    .B1(_08265_),
    .B2(_08271_),
    .X(_08272_));
 sky130_fd_sc_hd__a2bb2o_2 _22600_ (.A1_N(_08264_),
    .A2_N(_08272_),
    .B1(_08264_),
    .B2(_08272_),
    .X(_08273_));
 sky130_fd_sc_hd__a2bb2o_2 _22601_ (.A1_N(_08263_),
    .A2_N(_08273_),
    .B1(_08263_),
    .B2(_08273_),
    .X(_08274_));
 sky130_fd_sc_hd__a2bb2o_2 _22602_ (.A1_N(_08262_),
    .A2_N(_08274_),
    .B1(_08262_),
    .B2(_08274_),
    .X(_08275_));
 sky130_fd_sc_hd__o22a_2 _22603_ (.A1(_08140_),
    .A2(_08151_),
    .B1(_08139_),
    .B2(_08152_),
    .X(_08276_));
 sky130_fd_sc_hd__a2bb2o_2 _22604_ (.A1_N(_08275_),
    .A2_N(_08276_),
    .B1(_08275_),
    .B2(_08276_),
    .X(_08277_));
 sky130_fd_sc_hd__a2bb2o_2 _22605_ (.A1_N(_08261_),
    .A2_N(_08277_),
    .B1(_08261_),
    .B2(_08277_),
    .X(_08278_));
 sky130_fd_sc_hd__a2bb2o_2 _22606_ (.A1_N(_08258_),
    .A2_N(_08278_),
    .B1(_08258_),
    .B2(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__a2bb2o_2 _22607_ (.A1_N(_08257_),
    .A2_N(_08279_),
    .B1(_08257_),
    .B2(_08279_),
    .X(_08280_));
 sky130_fd_sc_hd__o22a_2 _22608_ (.A1(_08183_),
    .A2(_08184_),
    .B1(_08173_),
    .B2(_08185_),
    .X(_08281_));
 sky130_fd_sc_hd__o22a_2 _22609_ (.A1(_08190_),
    .A2(_08203_),
    .B1(_08189_),
    .B2(_08204_),
    .X(_08282_));
 sky130_fd_sc_hd__o22a_2 _22610_ (.A1(_08038_),
    .A2(_07007_),
    .B1(_04951_),
    .B2(_07009_),
    .X(_08283_));
 sky130_fd_sc_hd__and4_2 _22611_ (.A(_11614_),
    .B(_11882_),
    .C(_11617_),
    .D(_11880_),
    .X(_08284_));
 sky130_fd_sc_hd__nor2_2 _22612_ (.A(_08283_),
    .B(_08284_),
    .Y(_08285_));
 sky130_fd_sc_hd__nor2_2 _22613_ (.A(_04903_),
    .B(_07024_),
    .Y(_08286_));
 sky130_fd_sc_hd__a2bb2o_2 _22614_ (.A1_N(_08285_),
    .A2_N(_08286_),
    .B1(_08285_),
    .B2(_08286_),
    .X(_08287_));
 sky130_fd_sc_hd__or2_2 _22615_ (.A(_05133_),
    .B(_06878_),
    .X(_08288_));
 sky130_fd_sc_hd__o22a_2 _22616_ (.A1(_05945_),
    .A2(_06375_),
    .B1(_06415_),
    .B2(_06495_),
    .X(_08289_));
 sky130_fd_sc_hd__and4_2 _22617_ (.A(_06928_),
    .B(\pcpi_mul.rs1[25] ),
    .C(_06929_),
    .D(\pcpi_mul.rs1[26] ),
    .X(_08290_));
 sky130_fd_sc_hd__or2_2 _22618_ (.A(_08289_),
    .B(_08290_),
    .X(_08291_));
 sky130_fd_sc_hd__a2bb2o_2 _22619_ (.A1_N(_08288_),
    .A2_N(_08291_),
    .B1(_08288_),
    .B2(_08291_),
    .X(_08292_));
 sky130_fd_sc_hd__o21ba_2 _22620_ (.A1(_08166_),
    .A2(_08169_),
    .B1_N(_08168_),
    .X(_08293_));
 sky130_fd_sc_hd__a2bb2o_2 _22621_ (.A1_N(_08292_),
    .A2_N(_08293_),
    .B1(_08292_),
    .B2(_08293_),
    .X(_08294_));
 sky130_fd_sc_hd__a2bb2o_2 _22622_ (.A1_N(_08287_),
    .A2_N(_08294_),
    .B1(_08287_),
    .B2(_08294_),
    .X(_08295_));
 sky130_fd_sc_hd__a21oi_2 _22623_ (.A1(_08179_),
    .A2(_08180_),
    .B1(_08178_),
    .Y(_08296_));
 sky130_fd_sc_hd__o21ba_2 _22624_ (.A1(_08191_),
    .A2(_08194_),
    .B1_N(_08193_),
    .X(_08297_));
 sky130_fd_sc_hd__buf_1 _22625_ (.A(_06318_),
    .X(_08298_));
 sky130_fd_sc_hd__o22a_2 _22626_ (.A1(_08298_),
    .A2(_06904_),
    .B1(_08176_),
    .B2(_06754_),
    .X(_08299_));
 sky130_fd_sc_hd__buf_1 _22627_ (.A(_11602_),
    .X(_08300_));
 sky130_fd_sc_hd__buf_1 _22628_ (.A(_11605_),
    .X(_08301_));
 sky130_fd_sc_hd__and4_2 _22629_ (.A(_08300_),
    .B(_06499_),
    .C(_08301_),
    .D(_06627_),
    .X(_08302_));
 sky130_fd_sc_hd__nor2_2 _22630_ (.A(_08299_),
    .B(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__nor2_2 _22631_ (.A(_07922_),
    .B(_06234_),
    .Y(_08304_));
 sky130_fd_sc_hd__a2bb2o_2 _22632_ (.A1_N(_08303_),
    .A2_N(_08304_),
    .B1(_08303_),
    .B2(_08304_),
    .X(_08305_));
 sky130_fd_sc_hd__a2bb2o_2 _22633_ (.A1_N(_08297_),
    .A2_N(_08305_),
    .B1(_08297_),
    .B2(_08305_),
    .X(_08306_));
 sky130_fd_sc_hd__a2bb2o_2 _22634_ (.A1_N(_08296_),
    .A2_N(_08306_),
    .B1(_08296_),
    .B2(_08306_),
    .X(_08307_));
 sky130_fd_sc_hd__o22a_2 _22635_ (.A1(_08175_),
    .A2(_08181_),
    .B1(_08174_),
    .B2(_08182_),
    .X(_08308_));
 sky130_fd_sc_hd__a2bb2o_2 _22636_ (.A1_N(_08307_),
    .A2_N(_08308_),
    .B1(_08307_),
    .B2(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__a2bb2o_2 _22637_ (.A1_N(_08295_),
    .A2_N(_08309_),
    .B1(_08295_),
    .B2(_08309_),
    .X(_08310_));
 sky130_fd_sc_hd__a2bb2o_2 _22638_ (.A1_N(_08282_),
    .A2_N(_08310_),
    .B1(_08282_),
    .B2(_08310_),
    .X(_08311_));
 sky130_fd_sc_hd__a2bb2o_2 _22639_ (.A1_N(_08281_),
    .A2_N(_08311_),
    .B1(_08281_),
    .B2(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__o22a_2 _22640_ (.A1(_08200_),
    .A2(_08201_),
    .B1(_08195_),
    .B2(_08202_),
    .X(_08313_));
 sky130_fd_sc_hd__o22a_2 _22641_ (.A1(_08207_),
    .A2(_08212_),
    .B1(_08206_),
    .B2(_08213_),
    .X(_08314_));
 sky130_fd_sc_hd__or2_2 _22642_ (.A(_06700_),
    .B(_05987_),
    .X(_08315_));
 sky130_fd_sc_hd__o22a_2 _22643_ (.A1(_07359_),
    .A2(_05715_),
    .B1(_05662_),
    .B2(_05823_),
    .X(_08316_));
 sky130_fd_sc_hd__and4_2 _22644_ (.A(_06703_),
    .B(_06517_),
    .C(_06570_),
    .D(_06239_),
    .X(_08317_));
 sky130_fd_sc_hd__or2_2 _22645_ (.A(_08316_),
    .B(_08317_),
    .X(_08318_));
 sky130_fd_sc_hd__a2bb2o_2 _22646_ (.A1_N(_08315_),
    .A2_N(_08318_),
    .B1(_08315_),
    .B2(_08318_),
    .X(_08319_));
 sky130_fd_sc_hd__or2_2 _22647_ (.A(_07656_),
    .B(_06255_),
    .X(_08320_));
 sky130_fd_sc_hd__o22a_2 _22648_ (.A1(_07658_),
    .A2(_05501_),
    .B1(_06030_),
    .B2(_06257_),
    .X(_08321_));
 sky130_fd_sc_hd__and4_2 _22649_ (.A(_07515_),
    .B(_06138_),
    .C(_07516_),
    .D(_06392_),
    .X(_08322_));
 sky130_fd_sc_hd__or2_2 _22650_ (.A(_08321_),
    .B(_08322_),
    .X(_08323_));
 sky130_fd_sc_hd__a2bb2o_2 _22651_ (.A1_N(_08320_),
    .A2_N(_08323_),
    .B1(_08320_),
    .B2(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__o21ba_2 _22652_ (.A1(_08196_),
    .A2(_08199_),
    .B1_N(_08198_),
    .X(_08325_));
 sky130_fd_sc_hd__a2bb2o_2 _22653_ (.A1_N(_08324_),
    .A2_N(_08325_),
    .B1(_08324_),
    .B2(_08325_),
    .X(_08326_));
 sky130_fd_sc_hd__a2bb2o_2 _22654_ (.A1_N(_08319_),
    .A2_N(_08326_),
    .B1(_08319_),
    .B2(_08326_),
    .X(_08327_));
 sky130_fd_sc_hd__a2bb2o_2 _22655_ (.A1_N(_08314_),
    .A2_N(_08327_),
    .B1(_08314_),
    .B2(_08327_),
    .X(_08328_));
 sky130_fd_sc_hd__a2bb2o_2 _22656_ (.A1_N(_08313_),
    .A2_N(_08328_),
    .B1(_08313_),
    .B2(_08328_),
    .X(_08329_));
 sky130_fd_sc_hd__o21ba_2 _22657_ (.A1(_08208_),
    .A2(_08211_),
    .B1_N(_08210_),
    .X(_08330_));
 sky130_fd_sc_hd__o21ba_2 _22658_ (.A1(_08215_),
    .A2(_08218_),
    .B1_N(_08217_),
    .X(_08331_));
 sky130_fd_sc_hd__o22a_2 _22659_ (.A1(_07814_),
    .A2(_05169_),
    .B1(_06445_),
    .B2(_05256_),
    .X(_08332_));
 sky130_fd_sc_hd__and4_2 _22660_ (.A(_07816_),
    .B(_11923_),
    .C(_07672_),
    .D(_07509_),
    .X(_08333_));
 sky130_fd_sc_hd__nor2_2 _22661_ (.A(_08332_),
    .B(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__nor2_2 _22662_ (.A(_06447_),
    .B(_05421_),
    .Y(_08335_));
 sky130_fd_sc_hd__a2bb2o_2 _22663_ (.A1_N(_08334_),
    .A2_N(_08335_),
    .B1(_08334_),
    .B2(_08335_),
    .X(_08336_));
 sky130_fd_sc_hd__a2bb2o_2 _22664_ (.A1_N(_08331_),
    .A2_N(_08336_),
    .B1(_08331_),
    .B2(_08336_),
    .X(_08337_));
 sky130_fd_sc_hd__a2bb2o_2 _22665_ (.A1_N(_08330_),
    .A2_N(_08337_),
    .B1(_08330_),
    .B2(_08337_),
    .X(_08338_));
 sky130_fd_sc_hd__or2_2 _22666_ (.A(_06686_),
    .B(_05158_),
    .X(_08339_));
 sky130_fd_sc_hd__o22a_2 _22667_ (.A1(_07535_),
    .A2(_06180_),
    .B1(_07536_),
    .B2(_05530_),
    .X(_08340_));
 sky130_fd_sc_hd__and4_2 _22668_ (.A(_07538_),
    .B(_06184_),
    .C(_07539_),
    .D(_05743_),
    .X(_08341_));
 sky130_fd_sc_hd__or2_2 _22669_ (.A(_08340_),
    .B(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__a2bb2o_2 _22670_ (.A1_N(_08339_),
    .A2_N(_08342_),
    .B1(_08339_),
    .B2(_08342_),
    .X(_08343_));
 sky130_fd_sc_hd__or2_2 _22671_ (.A(_07828_),
    .B(_05943_),
    .X(_08344_));
 sky130_fd_sc_hd__and4_2 _22672_ (.A(_07830_),
    .B(_05190_),
    .C(_11560_),
    .D(_05578_),
    .X(_08345_));
 sky130_fd_sc_hd__o22a_2 _22673_ (.A1(_07832_),
    .A2(_05577_),
    .B1(_07965_),
    .B2(_05086_),
    .X(_08346_));
 sky130_fd_sc_hd__or2_2 _22674_ (.A(_08345_),
    .B(_08346_),
    .X(_08347_));
 sky130_fd_sc_hd__a2bb2o_2 _22675_ (.A1_N(_08344_),
    .A2_N(_08347_),
    .B1(_08344_),
    .B2(_08347_),
    .X(_08348_));
 sky130_fd_sc_hd__o21ba_2 _22676_ (.A1(_08220_),
    .A2(_08223_),
    .B1_N(_08221_),
    .X(_08349_));
 sky130_fd_sc_hd__a2bb2o_2 _22677_ (.A1_N(_08348_),
    .A2_N(_08349_),
    .B1(_08348_),
    .B2(_08349_),
    .X(_08350_));
 sky130_fd_sc_hd__a2bb2o_2 _22678_ (.A1_N(_08343_),
    .A2_N(_08350_),
    .B1(_08343_),
    .B2(_08350_),
    .X(_08351_));
 sky130_fd_sc_hd__o22a_2 _22679_ (.A1(_08224_),
    .A2(_08225_),
    .B1(_08219_),
    .B2(_08226_),
    .X(_08352_));
 sky130_fd_sc_hd__a2bb2o_2 _22680_ (.A1_N(_08351_),
    .A2_N(_08352_),
    .B1(_08351_),
    .B2(_08352_),
    .X(_08353_));
 sky130_fd_sc_hd__a2bb2o_2 _22681_ (.A1_N(_08338_),
    .A2_N(_08353_),
    .B1(_08338_),
    .B2(_08353_),
    .X(_08354_));
 sky130_fd_sc_hd__o22a_2 _22682_ (.A1(_08227_),
    .A2(_08228_),
    .B1(_08214_),
    .B2(_08229_),
    .X(_08355_));
 sky130_fd_sc_hd__a2bb2o_2 _22683_ (.A1_N(_08354_),
    .A2_N(_08355_),
    .B1(_08354_),
    .B2(_08355_),
    .X(_08356_));
 sky130_fd_sc_hd__a2bb2o_2 _22684_ (.A1_N(_08329_),
    .A2_N(_08356_),
    .B1(_08329_),
    .B2(_08356_),
    .X(_08357_));
 sky130_fd_sc_hd__o22a_2 _22685_ (.A1(_08230_),
    .A2(_08231_),
    .B1(_08205_),
    .B2(_08232_),
    .X(_08358_));
 sky130_fd_sc_hd__a2bb2o_2 _22686_ (.A1_N(_08357_),
    .A2_N(_08358_),
    .B1(_08357_),
    .B2(_08358_),
    .X(_08359_));
 sky130_fd_sc_hd__a2bb2o_2 _22687_ (.A1_N(_08312_),
    .A2_N(_08359_),
    .B1(_08312_),
    .B2(_08359_),
    .X(_08360_));
 sky130_fd_sc_hd__o22a_2 _22688_ (.A1(_08233_),
    .A2(_08234_),
    .B1(_08188_),
    .B2(_08235_),
    .X(_08361_));
 sky130_fd_sc_hd__a2bb2o_2 _22689_ (.A1_N(_08360_),
    .A2_N(_08361_),
    .B1(_08360_),
    .B2(_08361_),
    .X(_08362_));
 sky130_fd_sc_hd__a2bb2o_2 _22690_ (.A1_N(_08280_),
    .A2_N(_08362_),
    .B1(_08280_),
    .B2(_08362_),
    .X(_08363_));
 sky130_fd_sc_hd__o22a_2 _22691_ (.A1(_08236_),
    .A2(_08237_),
    .B1(_08158_),
    .B2(_08238_),
    .X(_08364_));
 sky130_fd_sc_hd__a2bb2o_2 _22692_ (.A1_N(_08363_),
    .A2_N(_08364_),
    .B1(_08363_),
    .B2(_08364_),
    .X(_08365_));
 sky130_fd_sc_hd__a2bb2o_2 _22693_ (.A1_N(_08256_),
    .A2_N(_08365_),
    .B1(_08256_),
    .B2(_08365_),
    .X(_08366_));
 sky130_fd_sc_hd__o22a_2 _22694_ (.A1(_08239_),
    .A2(_08240_),
    .B1(_08132_),
    .B2(_08241_),
    .X(_08367_));
 sky130_fd_sc_hd__a2bb2o_2 _22695_ (.A1_N(_08366_),
    .A2_N(_08367_),
    .B1(_08366_),
    .B2(_08367_),
    .X(_08368_));
 sky130_fd_sc_hd__a2bb2o_2 _22696_ (.A1_N(_08131_),
    .A2_N(_08368_),
    .B1(_08131_),
    .B2(_08368_),
    .X(_08369_));
 sky130_fd_sc_hd__a2bb2o_2 _22697_ (.A1_N(_08251_),
    .A2_N(_08369_),
    .B1(_08251_),
    .B2(_08369_),
    .X(_08370_));
 sky130_fd_sc_hd__o21ai_2 _22698_ (.A1(_08248_),
    .A2(_08250_),
    .B1(_08247_),
    .Y(_08371_));
 sky130_fd_sc_hd__a2bb2o_2 _22699_ (.A1_N(_08370_),
    .A2_N(_08371_),
    .B1(_08370_),
    .B2(_08371_),
    .X(_02658_));
 sky130_fd_sc_hd__o22a_2 _22700_ (.A1(_08258_),
    .A2(_08278_),
    .B1(_08257_),
    .B2(_08279_),
    .X(_08372_));
 sky130_fd_sc_hd__o21a_2 _22701_ (.A1(_08002_),
    .A2(_08259_),
    .B1(_08253_),
    .X(_08373_));
 sky130_fd_sc_hd__buf_1 _22702_ (.A(_08373_),
    .X(_08374_));
 sky130_fd_sc_hd__buf_1 _22703_ (.A(_08374_),
    .X(_08375_));
 sky130_fd_sc_hd__or2_2 _22704_ (.A(_08372_),
    .B(_08374_),
    .X(_08376_));
 sky130_fd_sc_hd__a21bo_2 _22705_ (.A1(_08372_),
    .A2(_08375_),
    .B1_N(_08376_),
    .X(_08377_));
 sky130_fd_sc_hd__buf_1 _22706_ (.A(_08260_),
    .X(_08378_));
 sky130_fd_sc_hd__buf_1 _22707_ (.A(_08378_),
    .X(_08379_));
 sky130_fd_sc_hd__o22a_2 _22708_ (.A1(_08275_),
    .A2(_08276_),
    .B1(_08379_),
    .B2(_08277_),
    .X(_08380_));
 sky130_fd_sc_hd__o22a_2 _22709_ (.A1(_08282_),
    .A2(_08310_),
    .B1(_08281_),
    .B2(_08311_),
    .X(_08381_));
 sky130_fd_sc_hd__o22a_2 _22710_ (.A1(_08265_),
    .A2(_08271_),
    .B1(_08264_),
    .B2(_08272_),
    .X(_08382_));
 sky130_fd_sc_hd__o22a_2 _22711_ (.A1(_08292_),
    .A2(_08293_),
    .B1(_08287_),
    .B2(_08294_),
    .X(_08383_));
 sky130_fd_sc_hd__o32a_2 _22712_ (.A1(_07602_),
    .A2(_07583_),
    .A3(_08268_),
    .B1(_08148_),
    .B2(_08270_),
    .X(_08384_));
 sky130_fd_sc_hd__a21oi_2 _22713_ (.A1(_08285_),
    .A2(_08286_),
    .B1(_08284_),
    .Y(_08385_));
 sky130_fd_sc_hd__or2_2 _22714_ (.A(_10584_),
    .B(_04865_),
    .X(_08386_));
 sky130_fd_sc_hd__a32o_2 _22715_ (.A1(_07868_),
    .A2(_11618_),
    .A3(_08269_),
    .B1(_08268_),
    .B2(_08386_),
    .X(_08387_));
 sky130_fd_sc_hd__a2bb2o_2 _22716_ (.A1_N(_08147_),
    .A2_N(_08387_),
    .B1(_08147_),
    .B2(_08387_),
    .X(_08388_));
 sky130_fd_sc_hd__buf_1 _22717_ (.A(_08388_),
    .X(_08389_));
 sky130_fd_sc_hd__buf_1 _22718_ (.A(_08388_),
    .X(_08390_));
 sky130_fd_sc_hd__a2bb2o_2 _22719_ (.A1_N(_08385_),
    .A2_N(_08389_),
    .B1(_08385_),
    .B2(_08390_),
    .X(_08391_));
 sky130_fd_sc_hd__a2bb2o_2 _22720_ (.A1_N(_08384_),
    .A2_N(_08391_),
    .B1(_08384_),
    .B2(_08391_),
    .X(_08392_));
 sky130_fd_sc_hd__a2bb2o_2 _22721_ (.A1_N(_08383_),
    .A2_N(_08392_),
    .B1(_08383_),
    .B2(_08392_),
    .X(_08393_));
 sky130_fd_sc_hd__a2bb2o_2 _22722_ (.A1_N(_08382_),
    .A2_N(_08393_),
    .B1(_08382_),
    .B2(_08393_),
    .X(_08394_));
 sky130_fd_sc_hd__o22a_2 _22723_ (.A1(_08263_),
    .A2(_08273_),
    .B1(_08262_),
    .B2(_08274_),
    .X(_08395_));
 sky130_fd_sc_hd__o2bb2ai_2 _22724_ (.A1_N(_08394_),
    .A2_N(_08395_),
    .B1(_08394_),
    .B2(_08395_),
    .Y(_08396_));
 sky130_fd_sc_hd__a2bb2o_2 _22725_ (.A1_N(_08261_),
    .A2_N(_08396_),
    .B1(_08261_),
    .B2(_08396_),
    .X(_08397_));
 sky130_fd_sc_hd__a2bb2o_2 _22726_ (.A1_N(_08381_),
    .A2_N(_08397_),
    .B1(_08381_),
    .B2(_08397_),
    .X(_08398_));
 sky130_fd_sc_hd__a2bb2o_2 _22727_ (.A1_N(_08380_),
    .A2_N(_08398_),
    .B1(_08380_),
    .B2(_08398_),
    .X(_08399_));
 sky130_fd_sc_hd__o22a_2 _22728_ (.A1(_08307_),
    .A2(_08308_),
    .B1(_08295_),
    .B2(_08309_),
    .X(_08400_));
 sky130_fd_sc_hd__o22a_2 _22729_ (.A1(_08314_),
    .A2(_08327_),
    .B1(_08313_),
    .B2(_08328_),
    .X(_08401_));
 sky130_fd_sc_hd__o22a_2 _22730_ (.A1(_08038_),
    .A2(_06890_),
    .B1(_04951_),
    .B2(_07022_),
    .X(_08402_));
 sky130_fd_sc_hd__and4_2 _22731_ (.A(_11614_),
    .B(_07587_),
    .C(_11617_),
    .D(_11876_),
    .X(_08403_));
 sky130_fd_sc_hd__nor2_2 _22732_ (.A(_08402_),
    .B(_08403_),
    .Y(_08404_));
 sky130_fd_sc_hd__nor2_2 _22733_ (.A(_04903_),
    .B(_08266_),
    .Y(_08405_));
 sky130_fd_sc_hd__a2bb2o_2 _22734_ (.A1_N(_08404_),
    .A2_N(_08405_),
    .B1(_08404_),
    .B2(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__o22a_2 _22735_ (.A1(_06178_),
    .A2(_06742_),
    .B1(_06179_),
    .B2(_06878_),
    .X(_08407_));
 sky130_fd_sc_hd__and4_2 _22736_ (.A(_07483_),
    .B(_07459_),
    .C(_07484_),
    .D(\pcpi_mul.rs1[27] ),
    .X(_08408_));
 sky130_fd_sc_hd__nor2_2 _22737_ (.A(_08407_),
    .B(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__nor2_2 _22738_ (.A(_06305_),
    .B(_07007_),
    .Y(_08410_));
 sky130_fd_sc_hd__a2bb2o_2 _22739_ (.A1_N(_08409_),
    .A2_N(_08410_),
    .B1(_08409_),
    .B2(_08410_),
    .X(_08411_));
 sky130_fd_sc_hd__o21ba_2 _22740_ (.A1(_08288_),
    .A2(_08291_),
    .B1_N(_08290_),
    .X(_08412_));
 sky130_fd_sc_hd__a2bb2o_2 _22741_ (.A1_N(_08411_),
    .A2_N(_08412_),
    .B1(_08411_),
    .B2(_08412_),
    .X(_08413_));
 sky130_fd_sc_hd__a2bb2o_2 _22742_ (.A1_N(_08406_),
    .A2_N(_08413_),
    .B1(_08406_),
    .B2(_08413_),
    .X(_08414_));
 sky130_fd_sc_hd__a21oi_2 _22743_ (.A1(_08303_),
    .A2(_08304_),
    .B1(_08302_),
    .Y(_08415_));
 sky130_fd_sc_hd__o21ba_2 _22744_ (.A1(_08315_),
    .A2(_08318_),
    .B1_N(_08317_),
    .X(_08416_));
 sky130_fd_sc_hd__o22a_2 _22745_ (.A1(_08298_),
    .A2(_06754_),
    .B1(_08176_),
    .B2(_06233_),
    .X(_08417_));
 sky130_fd_sc_hd__and4_2 _22746_ (.A(_08300_),
    .B(_06627_),
    .C(_08301_),
    .D(_06752_),
    .X(_08418_));
 sky130_fd_sc_hd__nor2_2 _22747_ (.A(_08417_),
    .B(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__nor2_2 _22748_ (.A(_07922_),
    .B(_06617_),
    .Y(_08420_));
 sky130_fd_sc_hd__a2bb2o_2 _22749_ (.A1_N(_08419_),
    .A2_N(_08420_),
    .B1(_08419_),
    .B2(_08420_),
    .X(_08421_));
 sky130_fd_sc_hd__a2bb2o_2 _22750_ (.A1_N(_08416_),
    .A2_N(_08421_),
    .B1(_08416_),
    .B2(_08421_),
    .X(_08422_));
 sky130_fd_sc_hd__a2bb2o_2 _22751_ (.A1_N(_08415_),
    .A2_N(_08422_),
    .B1(_08415_),
    .B2(_08422_),
    .X(_08423_));
 sky130_fd_sc_hd__o22a_2 _22752_ (.A1(_08297_),
    .A2(_08305_),
    .B1(_08296_),
    .B2(_08306_),
    .X(_08424_));
 sky130_fd_sc_hd__a2bb2o_2 _22753_ (.A1_N(_08423_),
    .A2_N(_08424_),
    .B1(_08423_),
    .B2(_08424_),
    .X(_08425_));
 sky130_fd_sc_hd__a2bb2o_2 _22754_ (.A1_N(_08414_),
    .A2_N(_08425_),
    .B1(_08414_),
    .B2(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__a2bb2o_2 _22755_ (.A1_N(_08401_),
    .A2_N(_08426_),
    .B1(_08401_),
    .B2(_08426_),
    .X(_08427_));
 sky130_fd_sc_hd__a2bb2o_2 _22756_ (.A1_N(_08400_),
    .A2_N(_08427_),
    .B1(_08400_),
    .B2(_08427_),
    .X(_08428_));
 sky130_fd_sc_hd__o22a_2 _22757_ (.A1(_08324_),
    .A2(_08325_),
    .B1(_08319_),
    .B2(_08326_),
    .X(_08429_));
 sky130_fd_sc_hd__o22a_2 _22758_ (.A1(_08331_),
    .A2(_08336_),
    .B1(_08330_),
    .B2(_08337_),
    .X(_08430_));
 sky130_fd_sc_hd__buf_1 _22759_ (.A(_05662_),
    .X(_08431_));
 sky130_fd_sc_hd__o22a_2 _22760_ (.A1(_07651_),
    .A2(_05884_),
    .B1(_08431_),
    .B2(_05892_),
    .X(_08432_));
 sky130_fd_sc_hd__buf_1 _22761_ (.A(_06703_),
    .X(_08433_));
 sky130_fd_sc_hd__buf_1 _22762_ (.A(_06570_),
    .X(_08434_));
 sky130_fd_sc_hd__and4_2 _22763_ (.A(_08433_),
    .B(_06240_),
    .C(_08434_),
    .D(_06372_),
    .X(_08435_));
 sky130_fd_sc_hd__nor2_2 _22764_ (.A(_08432_),
    .B(_08435_),
    .Y(_08436_));
 sky130_fd_sc_hd__buf_1 _22765_ (.A(_06700_),
    .X(_08437_));
 sky130_fd_sc_hd__nor2_2 _22766_ (.A(_08437_),
    .B(_08057_),
    .Y(_08438_));
 sky130_fd_sc_hd__a2bb2o_2 _22767_ (.A1_N(_08436_),
    .A2_N(_08438_),
    .B1(_08436_),
    .B2(_08438_),
    .X(_08439_));
 sky130_fd_sc_hd__buf_1 _22768_ (.A(_06579_),
    .X(_08440_));
 sky130_fd_sc_hd__buf_1 _22769_ (.A(_06033_),
    .X(_08441_));
 sky130_fd_sc_hd__o22a_2 _22770_ (.A1(_08440_),
    .A2(_05598_),
    .B1(_08441_),
    .B2(_07059_),
    .X(_08442_));
 sky130_fd_sc_hd__and4_2 _22771_ (.A(_07801_),
    .B(_05897_),
    .C(_07802_),
    .D(_05999_),
    .X(_08443_));
 sky130_fd_sc_hd__nor2_2 _22772_ (.A(_08442_),
    .B(_08443_),
    .Y(_08444_));
 sky130_fd_sc_hd__buf_1 _22773_ (.A(_06035_),
    .X(_08445_));
 sky130_fd_sc_hd__nor2_2 _22774_ (.A(_08445_),
    .B(_05716_),
    .Y(_08446_));
 sky130_fd_sc_hd__a2bb2o_2 _22775_ (.A1_N(_08444_),
    .A2_N(_08446_),
    .B1(_08444_),
    .B2(_08446_),
    .X(_08447_));
 sky130_fd_sc_hd__o21ba_2 _22776_ (.A1(_08320_),
    .A2(_08323_),
    .B1_N(_08322_),
    .X(_08448_));
 sky130_fd_sc_hd__a2bb2o_2 _22777_ (.A1_N(_08447_),
    .A2_N(_08448_),
    .B1(_08447_),
    .B2(_08448_),
    .X(_08449_));
 sky130_fd_sc_hd__a2bb2o_2 _22778_ (.A1_N(_08439_),
    .A2_N(_08449_),
    .B1(_08439_),
    .B2(_08449_),
    .X(_08450_));
 sky130_fd_sc_hd__a2bb2o_2 _22779_ (.A1_N(_08430_),
    .A2_N(_08450_),
    .B1(_08430_),
    .B2(_08450_),
    .X(_08451_));
 sky130_fd_sc_hd__a2bb2o_2 _22780_ (.A1_N(_08429_),
    .A2_N(_08451_),
    .B1(_08429_),
    .B2(_08451_),
    .X(_08452_));
 sky130_fd_sc_hd__a21oi_2 _22781_ (.A1(_08334_),
    .A2(_08335_),
    .B1(_08333_),
    .Y(_08453_));
 sky130_fd_sc_hd__o21ba_2 _22782_ (.A1(_08339_),
    .A2(_08342_),
    .B1_N(_08341_),
    .X(_08454_));
 sky130_fd_sc_hd__o22a_2 _22783_ (.A1(_07814_),
    .A2(_05256_),
    .B1(_06442_),
    .B2(_05343_),
    .X(_08455_));
 sky130_fd_sc_hd__buf_1 _22784_ (.A(_11580_),
    .X(_08456_));
 sky130_fd_sc_hd__and4_2 _22785_ (.A(_11575_),
    .B(_07509_),
    .C(_08456_),
    .D(_05830_),
    .X(_08457_));
 sky130_fd_sc_hd__nor2_2 _22786_ (.A(_08455_),
    .B(_08457_),
    .Y(_08458_));
 sky130_fd_sc_hd__nor2_2 _22787_ (.A(_06273_),
    .B(_05502_),
    .Y(_08459_));
 sky130_fd_sc_hd__a2bb2o_2 _22788_ (.A1_N(_08458_),
    .A2_N(_08459_),
    .B1(_08458_),
    .B2(_08459_),
    .X(_08460_));
 sky130_fd_sc_hd__a2bb2o_2 _22789_ (.A1_N(_08454_),
    .A2_N(_08460_),
    .B1(_08454_),
    .B2(_08460_),
    .X(_08461_));
 sky130_fd_sc_hd__a2bb2o_2 _22790_ (.A1_N(_08453_),
    .A2_N(_08461_),
    .B1(_08453_),
    .B2(_08461_),
    .X(_08462_));
 sky130_fd_sc_hd__or2_2 _22791_ (.A(_06686_),
    .B(_05736_),
    .X(_08463_));
 sky130_fd_sc_hd__o22a_2 _22792_ (.A1(_07535_),
    .A2(_05154_),
    .B1(_07536_),
    .B2(_05740_),
    .X(_08464_));
 sky130_fd_sc_hd__and4_2 _22793_ (.A(_07538_),
    .B(_05433_),
    .C(_07539_),
    .D(_05514_),
    .X(_08465_));
 sky130_fd_sc_hd__or2_2 _22794_ (.A(_08464_),
    .B(_08465_),
    .X(_08466_));
 sky130_fd_sc_hd__a2bb2o_2 _22795_ (.A1_N(_08463_),
    .A2_N(_08466_),
    .B1(_08463_),
    .B2(_08466_),
    .X(_08467_));
 sky130_fd_sc_hd__or2_2 _22796_ (.A(_07828_),
    .B(_05070_),
    .X(_08468_));
 sky130_fd_sc_hd__and4_2 _22797_ (.A(_07830_),
    .B(_05086_),
    .C(_08100_),
    .D(_11930_),
    .X(_08469_));
 sky130_fd_sc_hd__o22a_2 _22798_ (.A1(_07832_),
    .A2(_05578_),
    .B1(_07965_),
    .B2(_05076_),
    .X(_08470_));
 sky130_fd_sc_hd__or2_2 _22799_ (.A(_08469_),
    .B(_08470_),
    .X(_08471_));
 sky130_fd_sc_hd__a2bb2o_2 _22800_ (.A1_N(_08468_),
    .A2_N(_08471_),
    .B1(_08468_),
    .B2(_08471_),
    .X(_08472_));
 sky130_fd_sc_hd__o21ba_2 _22801_ (.A1(_08344_),
    .A2(_08347_),
    .B1_N(_08345_),
    .X(_08473_));
 sky130_fd_sc_hd__a2bb2o_2 _22802_ (.A1_N(_08472_),
    .A2_N(_08473_),
    .B1(_08472_),
    .B2(_08473_),
    .X(_08474_));
 sky130_fd_sc_hd__a2bb2o_2 _22803_ (.A1_N(_08467_),
    .A2_N(_08474_),
    .B1(_08467_),
    .B2(_08474_),
    .X(_08475_));
 sky130_fd_sc_hd__o22a_2 _22804_ (.A1(_08348_),
    .A2(_08349_),
    .B1(_08343_),
    .B2(_08350_),
    .X(_08476_));
 sky130_fd_sc_hd__a2bb2o_2 _22805_ (.A1_N(_08475_),
    .A2_N(_08476_),
    .B1(_08475_),
    .B2(_08476_),
    .X(_08477_));
 sky130_fd_sc_hd__a2bb2o_2 _22806_ (.A1_N(_08462_),
    .A2_N(_08477_),
    .B1(_08462_),
    .B2(_08477_),
    .X(_08478_));
 sky130_fd_sc_hd__o22a_2 _22807_ (.A1(_08351_),
    .A2(_08352_),
    .B1(_08338_),
    .B2(_08353_),
    .X(_08479_));
 sky130_fd_sc_hd__a2bb2o_2 _22808_ (.A1_N(_08478_),
    .A2_N(_08479_),
    .B1(_08478_),
    .B2(_08479_),
    .X(_08480_));
 sky130_fd_sc_hd__a2bb2o_2 _22809_ (.A1_N(_08452_),
    .A2_N(_08480_),
    .B1(_08452_),
    .B2(_08480_),
    .X(_08481_));
 sky130_fd_sc_hd__o22a_2 _22810_ (.A1(_08354_),
    .A2(_08355_),
    .B1(_08329_),
    .B2(_08356_),
    .X(_08482_));
 sky130_fd_sc_hd__a2bb2o_2 _22811_ (.A1_N(_08481_),
    .A2_N(_08482_),
    .B1(_08481_),
    .B2(_08482_),
    .X(_08483_));
 sky130_fd_sc_hd__a2bb2o_2 _22812_ (.A1_N(_08428_),
    .A2_N(_08483_),
    .B1(_08428_),
    .B2(_08483_),
    .X(_08484_));
 sky130_fd_sc_hd__o22a_2 _22813_ (.A1(_08357_),
    .A2(_08358_),
    .B1(_08312_),
    .B2(_08359_),
    .X(_08485_));
 sky130_fd_sc_hd__a2bb2o_2 _22814_ (.A1_N(_08484_),
    .A2_N(_08485_),
    .B1(_08484_),
    .B2(_08485_),
    .X(_08486_));
 sky130_fd_sc_hd__a2bb2o_2 _22815_ (.A1_N(_08399_),
    .A2_N(_08486_),
    .B1(_08399_),
    .B2(_08486_),
    .X(_08487_));
 sky130_fd_sc_hd__o22a_2 _22816_ (.A1(_08360_),
    .A2(_08361_),
    .B1(_08280_),
    .B2(_08362_),
    .X(_08488_));
 sky130_fd_sc_hd__a2bb2o_2 _22817_ (.A1_N(_08487_),
    .A2_N(_08488_),
    .B1(_08487_),
    .B2(_08488_),
    .X(_08489_));
 sky130_fd_sc_hd__a2bb2o_2 _22818_ (.A1_N(_08377_),
    .A2_N(_08489_),
    .B1(_08377_),
    .B2(_08489_),
    .X(_08490_));
 sky130_fd_sc_hd__o22a_2 _22819_ (.A1(_08363_),
    .A2(_08364_),
    .B1(_08256_),
    .B2(_08365_),
    .X(_08491_));
 sky130_fd_sc_hd__a2bb2o_2 _22820_ (.A1_N(_08490_),
    .A2_N(_08491_),
    .B1(_08490_),
    .B2(_08491_),
    .X(_08492_));
 sky130_fd_sc_hd__a2bb2o_2 _22821_ (.A1_N(_08255_),
    .A2_N(_08492_),
    .B1(_08255_),
    .B2(_08492_),
    .X(_08493_));
 sky130_fd_sc_hd__o22a_2 _22822_ (.A1(_08366_),
    .A2(_08367_),
    .B1(_08131_),
    .B2(_08368_),
    .X(_08494_));
 sky130_fd_sc_hd__or2_2 _22823_ (.A(_08493_),
    .B(_08494_),
    .X(_08495_));
 sky130_fd_sc_hd__a21bo_2 _22824_ (.A1(_08493_),
    .A2(_08494_),
    .B1_N(_08495_),
    .X(_08496_));
 sky130_fd_sc_hd__or2_2 _22825_ (.A(_08248_),
    .B(_08370_),
    .X(_08497_));
 sky130_fd_sc_hd__or3_2 _22826_ (.A(_07992_),
    .B(_08127_),
    .C(_08497_),
    .X(_08498_));
 sky130_fd_sc_hd__or2_2 _22827_ (.A(_07994_),
    .B(_08498_),
    .X(_08499_));
 sky130_fd_sc_hd__and2_2 _22828_ (.A(_08251_),
    .B(_08369_),
    .X(_08500_));
 sky130_fd_sc_hd__o22a_2 _22829_ (.A1(_08251_),
    .A2(_08369_),
    .B1(_08247_),
    .B2(_08500_),
    .X(_08501_));
 sky130_fd_sc_hd__o221a_2 _22830_ (.A1(_08249_),
    .A2(_08497_),
    .B1(_07996_),
    .B2(_08498_),
    .C1(_08501_),
    .X(_08502_));
 sky130_fd_sc_hd__o21ai_2 _22831_ (.A1(_07426_),
    .A2(_08499_),
    .B1(_08502_),
    .Y(_08503_));
 sky130_vsdinv _22832_ (.A(_08503_),
    .Y(_08504_));
 sky130_vsdinv _22833_ (.A(_08496_),
    .Y(_08505_));
 sky130_fd_sc_hd__o22a_2 _22834_ (.A1(_08496_),
    .A2(_08504_),
    .B1(_08505_),
    .B2(_08503_),
    .X(_02659_));
 sky130_fd_sc_hd__o22a_2 _22835_ (.A1(_08490_),
    .A2(_08491_),
    .B1(_08255_),
    .B2(_08492_),
    .X(_08506_));
 sky130_fd_sc_hd__o22a_2 _22836_ (.A1(_08381_),
    .A2(_08397_),
    .B1(_08380_),
    .B2(_08398_),
    .X(_08507_));
 sky130_fd_sc_hd__or2_2 _22837_ (.A(_08374_),
    .B(_08507_),
    .X(_08508_));
 sky130_fd_sc_hd__a21bo_2 _22838_ (.A1(_08375_),
    .A2(_08507_),
    .B1_N(_08508_),
    .X(_08509_));
 sky130_fd_sc_hd__o22a_2 _22839_ (.A1(_08394_),
    .A2(_08395_),
    .B1(_08379_),
    .B2(_08396_),
    .X(_08510_));
 sky130_fd_sc_hd__o22a_2 _22840_ (.A1(_08401_),
    .A2(_08426_),
    .B1(_08400_),
    .B2(_08427_),
    .X(_08511_));
 sky130_fd_sc_hd__buf_1 _22841_ (.A(_08260_),
    .X(_08512_));
 sky130_fd_sc_hd__o22a_2 _22842_ (.A1(_08385_),
    .A2(_08389_),
    .B1(_08384_),
    .B2(_08391_),
    .X(_08513_));
 sky130_fd_sc_hd__o22a_2 _22843_ (.A1(_08411_),
    .A2(_08412_),
    .B1(_08406_),
    .B2(_08413_),
    .X(_08514_));
 sky130_fd_sc_hd__o22a_2 _22844_ (.A1(_08268_),
    .A2(_08386_),
    .B1(_08148_),
    .B2(_08387_),
    .X(_08515_));
 sky130_fd_sc_hd__a21oi_2 _22845_ (.A1(_08404_),
    .A2(_08405_),
    .B1(_08403_),
    .Y(_08516_));
 sky130_fd_sc_hd__a2bb2o_2 _22846_ (.A1_N(_08390_),
    .A2_N(_08516_),
    .B1(_08388_),
    .B2(_08516_),
    .X(_08517_));
 sky130_fd_sc_hd__a2bb2o_2 _22847_ (.A1_N(_08515_),
    .A2_N(_08517_),
    .B1(_08515_),
    .B2(_08517_),
    .X(_08518_));
 sky130_fd_sc_hd__a2bb2o_2 _22848_ (.A1_N(_08514_),
    .A2_N(_08518_),
    .B1(_08514_),
    .B2(_08518_),
    .X(_08519_));
 sky130_fd_sc_hd__a2bb2o_2 _22849_ (.A1_N(_08513_),
    .A2_N(_08519_),
    .B1(_08513_),
    .B2(_08519_),
    .X(_08520_));
 sky130_fd_sc_hd__o22a_2 _22850_ (.A1(_08383_),
    .A2(_08392_),
    .B1(_08382_),
    .B2(_08393_),
    .X(_08521_));
 sky130_fd_sc_hd__o2bb2ai_2 _22851_ (.A1_N(_08520_),
    .A2_N(_08521_),
    .B1(_08520_),
    .B2(_08521_),
    .Y(_08522_));
 sky130_fd_sc_hd__a2bb2o_2 _22852_ (.A1_N(_08512_),
    .A2_N(_08522_),
    .B1(_08512_),
    .B2(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__a2bb2o_2 _22853_ (.A1_N(_08511_),
    .A2_N(_08523_),
    .B1(_08511_),
    .B2(_08523_),
    .X(_08524_));
 sky130_fd_sc_hd__a2bb2o_2 _22854_ (.A1_N(_08510_),
    .A2_N(_08524_),
    .B1(_08510_),
    .B2(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__o22a_2 _22855_ (.A1(_08423_),
    .A2(_08424_),
    .B1(_08414_),
    .B2(_08425_),
    .X(_08526_));
 sky130_fd_sc_hd__o22a_2 _22856_ (.A1(_08430_),
    .A2(_08450_),
    .B1(_08429_),
    .B2(_08451_),
    .X(_08527_));
 sky130_fd_sc_hd__o22a_2 _22857_ (.A1(_05060_),
    .A2(_07022_),
    .B1(_05667_),
    .B2(_07732_),
    .X(_08528_));
 sky130_fd_sc_hd__and4_2 _22858_ (.A(_05669_),
    .B(\pcpi_mul.rs1[30] ),
    .C(_05670_),
    .D(\pcpi_mul.rs1[31] ),
    .X(_08529_));
 sky130_fd_sc_hd__or2_2 _22859_ (.A(_08528_),
    .B(_08529_),
    .X(_08530_));
 sky130_vsdinv _22860_ (.A(_08530_),
    .Y(_08531_));
 sky130_fd_sc_hd__or2_2 _22861_ (.A(_10584_),
    .B(_04901_),
    .X(_08532_));
 sky130_fd_sc_hd__buf_1 _22862_ (.A(_08532_),
    .X(_08533_));
 sky130_fd_sc_hd__a32o_2 _22863_ (.A1(_07870_),
    .A2(\pcpi_mul.rs2[9] ),
    .A3(_08531_),
    .B1(_08530_),
    .B2(_08533_),
    .X(_08534_));
 sky130_fd_sc_hd__o22a_2 _22864_ (.A1(_06178_),
    .A2(_06623_),
    .B1(_07481_),
    .B2(_06749_),
    .X(_08535_));
 sky130_fd_sc_hd__and4_2 _22865_ (.A(_07483_),
    .B(\pcpi_mul.rs1[27] ),
    .C(_07484_),
    .D(_07749_),
    .X(_08536_));
 sky130_fd_sc_hd__nor2_2 _22866_ (.A(_08535_),
    .B(_08536_),
    .Y(_08537_));
 sky130_fd_sc_hd__nor2_2 _22867_ (.A(_07624_),
    .B(_07009_),
    .Y(_08538_));
 sky130_fd_sc_hd__a2bb2o_2 _22868_ (.A1_N(_08537_),
    .A2_N(_08538_),
    .B1(_08537_),
    .B2(_08538_),
    .X(_08539_));
 sky130_fd_sc_hd__a21oi_2 _22869_ (.A1(_08409_),
    .A2(_08410_),
    .B1(_08408_),
    .Y(_08540_));
 sky130_fd_sc_hd__a2bb2o_2 _22870_ (.A1_N(_08539_),
    .A2_N(_08540_),
    .B1(_08539_),
    .B2(_08540_),
    .X(_08541_));
 sky130_fd_sc_hd__a2bb2o_2 _22871_ (.A1_N(_08534_),
    .A2_N(_08541_),
    .B1(_08534_),
    .B2(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__a21oi_2 _22872_ (.A1(_08419_),
    .A2(_08420_),
    .B1(_08418_),
    .Y(_08543_));
 sky130_fd_sc_hd__a21oi_2 _22873_ (.A1(_08436_),
    .A2(_08438_),
    .B1(_08435_),
    .Y(_08544_));
 sky130_fd_sc_hd__o22a_2 _22874_ (.A1(_08298_),
    .A2(_06233_),
    .B1(_05392_),
    .B2(_06616_),
    .X(_08545_));
 sky130_fd_sc_hd__and4_2 _22875_ (.A(_08300_),
    .B(_06752_),
    .C(_08301_),
    .D(_06885_),
    .X(_08546_));
 sky130_fd_sc_hd__nor2_2 _22876_ (.A(_08545_),
    .B(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__nor2_2 _22877_ (.A(_07346_),
    .B(_06497_),
    .Y(_08548_));
 sky130_fd_sc_hd__a2bb2o_2 _22878_ (.A1_N(_08547_),
    .A2_N(_08548_),
    .B1(_08547_),
    .B2(_08548_),
    .X(_08549_));
 sky130_fd_sc_hd__a2bb2o_2 _22879_ (.A1_N(_08544_),
    .A2_N(_08549_),
    .B1(_08544_),
    .B2(_08549_),
    .X(_08550_));
 sky130_fd_sc_hd__a2bb2o_2 _22880_ (.A1_N(_08543_),
    .A2_N(_08550_),
    .B1(_08543_),
    .B2(_08550_),
    .X(_08551_));
 sky130_fd_sc_hd__o22a_2 _22881_ (.A1(_08416_),
    .A2(_08421_),
    .B1(_08415_),
    .B2(_08422_),
    .X(_08552_));
 sky130_fd_sc_hd__a2bb2o_2 _22882_ (.A1_N(_08551_),
    .A2_N(_08552_),
    .B1(_08551_),
    .B2(_08552_),
    .X(_08553_));
 sky130_fd_sc_hd__a2bb2o_2 _22883_ (.A1_N(_08542_),
    .A2_N(_08553_),
    .B1(_08542_),
    .B2(_08553_),
    .X(_08554_));
 sky130_fd_sc_hd__a2bb2o_2 _22884_ (.A1_N(_08527_),
    .A2_N(_08554_),
    .B1(_08527_),
    .B2(_08554_),
    .X(_08555_));
 sky130_fd_sc_hd__a2bb2o_2 _22885_ (.A1_N(_08526_),
    .A2_N(_08555_),
    .B1(_08526_),
    .B2(_08555_),
    .X(_08556_));
 sky130_fd_sc_hd__o22a_2 _22886_ (.A1(_08447_),
    .A2(_08448_),
    .B1(_08439_),
    .B2(_08449_),
    .X(_08557_));
 sky130_fd_sc_hd__o22a_2 _22887_ (.A1(_08454_),
    .A2(_08460_),
    .B1(_08453_),
    .B2(_08461_),
    .X(_08558_));
 sky130_fd_sc_hd__buf_1 _22888_ (.A(_07359_),
    .X(_08559_));
 sky130_fd_sc_hd__o22a_2 _22889_ (.A1(_08559_),
    .A2(_05892_),
    .B1(_08431_),
    .B2(_05996_),
    .X(_08560_));
 sky130_fd_sc_hd__and4_2 _22890_ (.A(_08433_),
    .B(_06372_),
    .C(_08434_),
    .D(_11900_),
    .X(_08561_));
 sky130_fd_sc_hd__nor2_2 _22891_ (.A(_08560_),
    .B(_08561_),
    .Y(_08562_));
 sky130_fd_sc_hd__nor2_2 _22892_ (.A(_08437_),
    .B(_06360_),
    .Y(_08563_));
 sky130_fd_sc_hd__a2bb2o_2 _22893_ (.A1_N(_08562_),
    .A2_N(_08563_),
    .B1(_08562_),
    .B2(_08563_),
    .X(_08564_));
 sky130_fd_sc_hd__o22a_2 _22894_ (.A1(_08440_),
    .A2(_07059_),
    .B1(_08441_),
    .B2(_07196_),
    .X(_08565_));
 sky130_fd_sc_hd__and4_2 _22895_ (.A(_07801_),
    .B(_05999_),
    .C(_07802_),
    .D(_06117_),
    .X(_08566_));
 sky130_fd_sc_hd__nor2_2 _22896_ (.A(_08565_),
    .B(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__nor2_2 _22897_ (.A(_08445_),
    .B(_05824_),
    .Y(_08568_));
 sky130_fd_sc_hd__a2bb2o_2 _22898_ (.A1_N(_08567_),
    .A2_N(_08568_),
    .B1(_08567_),
    .B2(_08568_),
    .X(_08569_));
 sky130_fd_sc_hd__a21oi_2 _22899_ (.A1(_08444_),
    .A2(_08446_),
    .B1(_08443_),
    .Y(_08570_));
 sky130_fd_sc_hd__a2bb2o_2 _22900_ (.A1_N(_08569_),
    .A2_N(_08570_),
    .B1(_08569_),
    .B2(_08570_),
    .X(_08571_));
 sky130_fd_sc_hd__a2bb2o_2 _22901_ (.A1_N(_08564_),
    .A2_N(_08571_),
    .B1(_08564_),
    .B2(_08571_),
    .X(_08572_));
 sky130_fd_sc_hd__a2bb2o_2 _22902_ (.A1_N(_08558_),
    .A2_N(_08572_),
    .B1(_08558_),
    .B2(_08572_),
    .X(_08573_));
 sky130_fd_sc_hd__a2bb2o_2 _22903_ (.A1_N(_08557_),
    .A2_N(_08573_),
    .B1(_08557_),
    .B2(_08573_),
    .X(_08574_));
 sky130_fd_sc_hd__a21oi_2 _22904_ (.A1(_08458_),
    .A2(_08459_),
    .B1(_08457_),
    .Y(_08575_));
 sky130_fd_sc_hd__o21ba_2 _22905_ (.A1(_08463_),
    .A2(_08466_),
    .B1_N(_08465_),
    .X(_08576_));
 sky130_fd_sc_hd__o22a_2 _22906_ (.A1(_07814_),
    .A2(_05343_),
    .B1(_06445_),
    .B2(_05429_),
    .X(_08577_));
 sky130_fd_sc_hd__and4_2 _22907_ (.A(_07816_),
    .B(_05830_),
    .C(_08456_),
    .D(_05831_),
    .X(_08578_));
 sky130_fd_sc_hd__nor2_2 _22908_ (.A(_08577_),
    .B(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__nor2_2 _22909_ (.A(_06447_),
    .B(_05599_),
    .Y(_08580_));
 sky130_fd_sc_hd__a2bb2o_2 _22910_ (.A1_N(_08579_),
    .A2_N(_08580_),
    .B1(_08579_),
    .B2(_08580_),
    .X(_08581_));
 sky130_fd_sc_hd__a2bb2o_2 _22911_ (.A1_N(_08576_),
    .A2_N(_08581_),
    .B1(_08576_),
    .B2(_08581_),
    .X(_08582_));
 sky130_fd_sc_hd__a2bb2o_2 _22912_ (.A1_N(_08575_),
    .A2_N(_08582_),
    .B1(_08575_),
    .B2(_08582_),
    .X(_08583_));
 sky130_fd_sc_hd__buf_1 _22913_ (.A(_07387_),
    .X(_08584_));
 sky130_fd_sc_hd__o22a_2 _22914_ (.A1(_08584_),
    .A2(_05937_),
    .B1(_06833_),
    .B2(_05736_),
    .X(_08585_));
 sky130_fd_sc_hd__and4_2 _22915_ (.A(_07680_),
    .B(_11925_),
    .C(_07681_),
    .D(_11923_),
    .X(_08586_));
 sky130_fd_sc_hd__nor2_2 _22916_ (.A(_08585_),
    .B(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__nor2_2 _22917_ (.A(_07822_),
    .B(_05335_),
    .Y(_08588_));
 sky130_fd_sc_hd__a2bb2o_2 _22918_ (.A1_N(_08587_),
    .A2_N(_08588_),
    .B1(_08587_),
    .B2(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__or2_2 _22919_ (.A(_08098_),
    .B(_05072_),
    .X(_08590_));
 sky130_fd_sc_hd__and4_2 _22920_ (.A(_07686_),
    .B(_05076_),
    .C(_08100_),
    .D(_11928_),
    .X(_08591_));
 sky130_fd_sc_hd__buf_1 _22921_ (.A(_10596_),
    .X(_08592_));
 sky130_fd_sc_hd__o22a_2 _22922_ (.A1(_08592_),
    .A2(_05177_),
    .B1(_07965_),
    .B2(_05163_),
    .X(_08593_));
 sky130_fd_sc_hd__or2_2 _22923_ (.A(_08591_),
    .B(_08593_),
    .X(_08594_));
 sky130_fd_sc_hd__a2bb2o_2 _22924_ (.A1_N(_08590_),
    .A2_N(_08594_),
    .B1(_08590_),
    .B2(_08594_),
    .X(_08595_));
 sky130_fd_sc_hd__o21ba_2 _22925_ (.A1(_08468_),
    .A2(_08471_),
    .B1_N(_08469_),
    .X(_08596_));
 sky130_fd_sc_hd__a2bb2o_2 _22926_ (.A1_N(_08595_),
    .A2_N(_08596_),
    .B1(_08595_),
    .B2(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__a2bb2o_2 _22927_ (.A1_N(_08589_),
    .A2_N(_08597_),
    .B1(_08589_),
    .B2(_08597_),
    .X(_08598_));
 sky130_fd_sc_hd__o22a_2 _22928_ (.A1(_08472_),
    .A2(_08473_),
    .B1(_08467_),
    .B2(_08474_),
    .X(_08599_));
 sky130_fd_sc_hd__a2bb2o_2 _22929_ (.A1_N(_08598_),
    .A2_N(_08599_),
    .B1(_08598_),
    .B2(_08599_),
    .X(_08600_));
 sky130_fd_sc_hd__a2bb2o_2 _22930_ (.A1_N(_08583_),
    .A2_N(_08600_),
    .B1(_08583_),
    .B2(_08600_),
    .X(_08601_));
 sky130_fd_sc_hd__o22a_2 _22931_ (.A1(_08475_),
    .A2(_08476_),
    .B1(_08462_),
    .B2(_08477_),
    .X(_08602_));
 sky130_fd_sc_hd__a2bb2o_2 _22932_ (.A1_N(_08601_),
    .A2_N(_08602_),
    .B1(_08601_),
    .B2(_08602_),
    .X(_08603_));
 sky130_fd_sc_hd__a2bb2o_2 _22933_ (.A1_N(_08574_),
    .A2_N(_08603_),
    .B1(_08574_),
    .B2(_08603_),
    .X(_08604_));
 sky130_fd_sc_hd__o22a_2 _22934_ (.A1(_08478_),
    .A2(_08479_),
    .B1(_08452_),
    .B2(_08480_),
    .X(_08605_));
 sky130_fd_sc_hd__a2bb2o_2 _22935_ (.A1_N(_08604_),
    .A2_N(_08605_),
    .B1(_08604_),
    .B2(_08605_),
    .X(_08606_));
 sky130_fd_sc_hd__a2bb2o_2 _22936_ (.A1_N(_08556_),
    .A2_N(_08606_),
    .B1(_08556_),
    .B2(_08606_),
    .X(_08607_));
 sky130_fd_sc_hd__o22a_2 _22937_ (.A1(_08481_),
    .A2(_08482_),
    .B1(_08428_),
    .B2(_08483_),
    .X(_08608_));
 sky130_fd_sc_hd__a2bb2o_2 _22938_ (.A1_N(_08607_),
    .A2_N(_08608_),
    .B1(_08607_),
    .B2(_08608_),
    .X(_08609_));
 sky130_fd_sc_hd__a2bb2o_2 _22939_ (.A1_N(_08525_),
    .A2_N(_08609_),
    .B1(_08525_),
    .B2(_08609_),
    .X(_08610_));
 sky130_fd_sc_hd__o22a_2 _22940_ (.A1(_08484_),
    .A2(_08485_),
    .B1(_08399_),
    .B2(_08486_),
    .X(_08611_));
 sky130_fd_sc_hd__a2bb2o_2 _22941_ (.A1_N(_08610_),
    .A2_N(_08611_),
    .B1(_08610_),
    .B2(_08611_),
    .X(_08612_));
 sky130_fd_sc_hd__a2bb2o_2 _22942_ (.A1_N(_08509_),
    .A2_N(_08612_),
    .B1(_08509_),
    .B2(_08612_),
    .X(_08613_));
 sky130_fd_sc_hd__o22a_2 _22943_ (.A1(_08487_),
    .A2(_08488_),
    .B1(_08377_),
    .B2(_08489_),
    .X(_08614_));
 sky130_fd_sc_hd__a2bb2o_2 _22944_ (.A1_N(_08613_),
    .A2_N(_08614_),
    .B1(_08613_),
    .B2(_08614_),
    .X(_08615_));
 sky130_fd_sc_hd__a2bb2o_2 _22945_ (.A1_N(_08376_),
    .A2_N(_08615_),
    .B1(_08376_),
    .B2(_08615_),
    .X(_08616_));
 sky130_fd_sc_hd__or2_2 _22946_ (.A(_08506_),
    .B(_08616_),
    .X(_08617_));
 sky130_fd_sc_hd__a21bo_2 _22947_ (.A1(_08506_),
    .A2(_08616_),
    .B1_N(_08617_),
    .X(_08618_));
 sky130_fd_sc_hd__o21ai_2 _22948_ (.A1(_08496_),
    .A2(_08504_),
    .B1(_08495_),
    .Y(_08619_));
 sky130_fd_sc_hd__a2bb2o_2 _22949_ (.A1_N(_08618_),
    .A2_N(_08619_),
    .B1(_08618_),
    .B2(_08619_),
    .X(_02660_));
 sky130_fd_sc_hd__o22a_2 _22950_ (.A1(_08511_),
    .A2(_08523_),
    .B1(_08510_),
    .B2(_08524_),
    .X(_08620_));
 sky130_fd_sc_hd__or2_2 _22951_ (.A(_08373_),
    .B(_08620_),
    .X(_08621_));
 sky130_fd_sc_hd__a21bo_2 _22952_ (.A1(_08375_),
    .A2(_08620_),
    .B1_N(_08621_),
    .X(_08622_));
 sky130_fd_sc_hd__buf_1 _22953_ (.A(_08260_),
    .X(_08623_));
 sky130_fd_sc_hd__o22a_2 _22954_ (.A1(_08520_),
    .A2(_08521_),
    .B1(_08623_),
    .B2(_08522_),
    .X(_08624_));
 sky130_fd_sc_hd__o22a_2 _22955_ (.A1(_08527_),
    .A2(_08554_),
    .B1(_08526_),
    .B2(_08555_),
    .X(_08625_));
 sky130_fd_sc_hd__o22a_2 _22956_ (.A1(_08539_),
    .A2(_08540_),
    .B1(_08534_),
    .B2(_08541_),
    .X(_08626_));
 sky130_fd_sc_hd__buf_1 _22957_ (.A(_08515_),
    .X(_08627_));
 sky130_fd_sc_hd__o21ba_2 _22958_ (.A1(_08530_),
    .A2(_08532_),
    .B1_N(_08529_),
    .X(_08628_));
 sky130_fd_sc_hd__a2bb2o_2 _22959_ (.A1_N(_08390_),
    .A2_N(_08628_),
    .B1(_08390_),
    .B2(_08628_),
    .X(_08629_));
 sky130_fd_sc_hd__a2bb2o_2 _22960_ (.A1_N(_08627_),
    .A2_N(_08629_),
    .B1(_08515_),
    .B2(_08629_),
    .X(_08630_));
 sky130_fd_sc_hd__o2bb2ai_2 _22961_ (.A1_N(_08626_),
    .A2_N(_08630_),
    .B1(_08626_),
    .B2(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__o22a_2 _22962_ (.A1(_08389_),
    .A2(_08516_),
    .B1(_08627_),
    .B2(_08517_),
    .X(_08632_));
 sky130_fd_sc_hd__o2bb2a_2 _22963_ (.A1_N(_08631_),
    .A2_N(_08632_),
    .B1(_08631_),
    .B2(_08632_),
    .X(_08633_));
 sky130_vsdinv _22964_ (.A(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__o22a_2 _22965_ (.A1(_08514_),
    .A2(_08518_),
    .B1(_08513_),
    .B2(_08519_),
    .X(_08635_));
 sky130_vsdinv _22966_ (.A(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__a22o_2 _22967_ (.A1(_08634_),
    .A2(_08635_),
    .B1(_08633_),
    .B2(_08636_),
    .X(_08637_));
 sky130_fd_sc_hd__a2bb2o_2 _22968_ (.A1_N(_08378_),
    .A2_N(_08637_),
    .B1(_08378_),
    .B2(_08637_),
    .X(_08638_));
 sky130_fd_sc_hd__a2bb2o_2 _22969_ (.A1_N(_08625_),
    .A2_N(_08638_),
    .B1(_08625_),
    .B2(_08638_),
    .X(_08639_));
 sky130_fd_sc_hd__a2bb2o_2 _22970_ (.A1_N(_08624_),
    .A2_N(_08639_),
    .B1(_08624_),
    .B2(_08639_),
    .X(_08640_));
 sky130_fd_sc_hd__o22a_2 _22971_ (.A1(_08551_),
    .A2(_08552_),
    .B1(_08542_),
    .B2(_08553_),
    .X(_08641_));
 sky130_fd_sc_hd__o22a_2 _22972_ (.A1(_08558_),
    .A2(_08572_),
    .B1(_08557_),
    .B2(_08573_),
    .X(_08642_));
 sky130_fd_sc_hd__nor2_2 _22973_ (.A(_08038_),
    .B(_07159_),
    .Y(_08643_));
 sky130_fd_sc_hd__or2_2 _22974_ (.A(_10584_),
    .B(_04949_),
    .X(_08644_));
 sky130_vsdinv _22975_ (.A(_08644_),
    .Y(_08645_));
 sky130_fd_sc_hd__a2bb2o_2 _22976_ (.A1_N(_08643_),
    .A2_N(_08645_),
    .B1(_08643_),
    .B2(_08645_),
    .X(_08646_));
 sky130_fd_sc_hd__a2bb2o_2 _22977_ (.A1_N(_08533_),
    .A2_N(_08646_),
    .B1(_08533_),
    .B2(_08646_),
    .X(_08647_));
 sky130_fd_sc_hd__o22a_2 _22978_ (.A1(_06178_),
    .A2(_06748_),
    .B1(_07481_),
    .B2(_06890_),
    .X(_08648_));
 sky130_fd_sc_hd__and4_2 _22979_ (.A(_07483_),
    .B(_07749_),
    .C(_07484_),
    .D(_07587_),
    .X(_08649_));
 sky130_fd_sc_hd__nor2_2 _22980_ (.A(_08648_),
    .B(_08649_),
    .Y(_08650_));
 sky130_fd_sc_hd__nor2_2 _22981_ (.A(_07624_),
    .B(_07023_),
    .Y(_08651_));
 sky130_fd_sc_hd__a2bb2o_2 _22982_ (.A1_N(_08650_),
    .A2_N(_08651_),
    .B1(_08650_),
    .B2(_08651_),
    .X(_08652_));
 sky130_fd_sc_hd__a21oi_2 _22983_ (.A1(_08537_),
    .A2(_08538_),
    .B1(_08536_),
    .Y(_08653_));
 sky130_fd_sc_hd__a2bb2o_2 _22984_ (.A1_N(_08652_),
    .A2_N(_08653_),
    .B1(_08652_),
    .B2(_08653_),
    .X(_08654_));
 sky130_fd_sc_hd__a2bb2o_2 _22985_ (.A1_N(_08647_),
    .A2_N(_08654_),
    .B1(_08647_),
    .B2(_08654_),
    .X(_08655_));
 sky130_fd_sc_hd__a21oi_2 _22986_ (.A1(_08547_),
    .A2(_08548_),
    .B1(_08546_),
    .Y(_08656_));
 sky130_fd_sc_hd__a21oi_2 _22987_ (.A1(_08562_),
    .A2(_08563_),
    .B1(_08561_),
    .Y(_08657_));
 sky130_fd_sc_hd__o22a_2 _22988_ (.A1(_08298_),
    .A2(_06616_),
    .B1(_08176_),
    .B2(_06496_),
    .X(_08658_));
 sky130_fd_sc_hd__and4_2 _22989_ (.A(_08300_),
    .B(_06885_),
    .C(_08301_),
    .D(_07459_),
    .X(_08659_));
 sky130_fd_sc_hd__nor2_2 _22990_ (.A(_08658_),
    .B(_08659_),
    .Y(_08660_));
 sky130_fd_sc_hd__nor2_2 _22991_ (.A(_07922_),
    .B(_06625_),
    .Y(_08661_));
 sky130_fd_sc_hd__a2bb2o_2 _22992_ (.A1_N(_08660_),
    .A2_N(_08661_),
    .B1(_08660_),
    .B2(_08661_),
    .X(_08662_));
 sky130_fd_sc_hd__a2bb2o_2 _22993_ (.A1_N(_08657_),
    .A2_N(_08662_),
    .B1(_08657_),
    .B2(_08662_),
    .X(_08663_));
 sky130_fd_sc_hd__a2bb2o_2 _22994_ (.A1_N(_08656_),
    .A2_N(_08663_),
    .B1(_08656_),
    .B2(_08663_),
    .X(_08664_));
 sky130_fd_sc_hd__o22a_2 _22995_ (.A1(_08544_),
    .A2(_08549_),
    .B1(_08543_),
    .B2(_08550_),
    .X(_08665_));
 sky130_fd_sc_hd__a2bb2o_2 _22996_ (.A1_N(_08664_),
    .A2_N(_08665_),
    .B1(_08664_),
    .B2(_08665_),
    .X(_08666_));
 sky130_fd_sc_hd__a2bb2o_2 _22997_ (.A1_N(_08655_),
    .A2_N(_08666_),
    .B1(_08655_),
    .B2(_08666_),
    .X(_08667_));
 sky130_fd_sc_hd__a2bb2o_2 _22998_ (.A1_N(_08642_),
    .A2_N(_08667_),
    .B1(_08642_),
    .B2(_08667_),
    .X(_08668_));
 sky130_fd_sc_hd__a2bb2o_2 _22999_ (.A1_N(_08641_),
    .A2_N(_08668_),
    .B1(_08641_),
    .B2(_08668_),
    .X(_08669_));
 sky130_fd_sc_hd__o22a_2 _23000_ (.A1(_08569_),
    .A2(_08570_),
    .B1(_08564_),
    .B2(_08571_),
    .X(_08670_));
 sky130_fd_sc_hd__o22a_2 _23001_ (.A1(_08576_),
    .A2(_08581_),
    .B1(_08575_),
    .B2(_08582_),
    .X(_08671_));
 sky130_fd_sc_hd__o22a_2 _23002_ (.A1(_08559_),
    .A2(_06502_),
    .B1(_08431_),
    .B2(_06359_),
    .X(_08672_));
 sky130_fd_sc_hd__and4_2 _23003_ (.A(_08433_),
    .B(_11900_),
    .C(_08434_),
    .D(_11897_),
    .X(_08673_));
 sky130_fd_sc_hd__nor2_2 _23004_ (.A(_08672_),
    .B(_08673_),
    .Y(_08674_));
 sky130_fd_sc_hd__nor2_2 _23005_ (.A(_08437_),
    .B(_06362_),
    .Y(_08675_));
 sky130_fd_sc_hd__a2bb2o_2 _23006_ (.A1_N(_08674_),
    .A2_N(_08675_),
    .B1(_08674_),
    .B2(_08675_),
    .X(_08676_));
 sky130_fd_sc_hd__o22a_2 _23007_ (.A1(_08440_),
    .A2(_07196_),
    .B1(_08441_),
    .B2(_05823_),
    .X(_08677_));
 sky130_fd_sc_hd__and4_2 _23008_ (.A(_07801_),
    .B(_11908_),
    .C(_07802_),
    .D(_11905_),
    .X(_08678_));
 sky130_fd_sc_hd__nor2_2 _23009_ (.A(_08677_),
    .B(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__nor2_2 _23010_ (.A(_08445_),
    .B(_05893_),
    .Y(_08680_));
 sky130_fd_sc_hd__a2bb2o_2 _23011_ (.A1_N(_08679_),
    .A2_N(_08680_),
    .B1(_08679_),
    .B2(_08680_),
    .X(_08681_));
 sky130_fd_sc_hd__a21oi_2 _23012_ (.A1(_08567_),
    .A2(_08568_),
    .B1(_08566_),
    .Y(_08682_));
 sky130_fd_sc_hd__a2bb2o_2 _23013_ (.A1_N(_08681_),
    .A2_N(_08682_),
    .B1(_08681_),
    .B2(_08682_),
    .X(_08683_));
 sky130_fd_sc_hd__a2bb2o_2 _23014_ (.A1_N(_08676_),
    .A2_N(_08683_),
    .B1(_08676_),
    .B2(_08683_),
    .X(_08684_));
 sky130_fd_sc_hd__a2bb2o_2 _23015_ (.A1_N(_08671_),
    .A2_N(_08684_),
    .B1(_08671_),
    .B2(_08684_),
    .X(_08685_));
 sky130_fd_sc_hd__a2bb2o_2 _23016_ (.A1_N(_08670_),
    .A2_N(_08685_),
    .B1(_08670_),
    .B2(_08685_),
    .X(_08686_));
 sky130_fd_sc_hd__a21oi_2 _23017_ (.A1(_08579_),
    .A2(_08580_),
    .B1(_08578_),
    .Y(_08687_));
 sky130_fd_sc_hd__a21oi_2 _23018_ (.A1(_08587_),
    .A2(_08588_),
    .B1(_08586_),
    .Y(_08688_));
 sky130_fd_sc_hd__o22a_2 _23019_ (.A1(_07814_),
    .A2(_06134_),
    .B1(_06445_),
    .B2(_05895_),
    .X(_08689_));
 sky130_fd_sc_hd__and4_2 _23020_ (.A(_07816_),
    .B(_05831_),
    .C(_08456_),
    .D(_05897_),
    .X(_08690_));
 sky130_fd_sc_hd__nor2_2 _23021_ (.A(_08689_),
    .B(_08690_),
    .Y(_08691_));
 sky130_fd_sc_hd__nor2_2 _23022_ (.A(_06447_),
    .B(_05704_),
    .Y(_08692_));
 sky130_fd_sc_hd__a2bb2o_2 _23023_ (.A1_N(_08691_),
    .A2_N(_08692_),
    .B1(_08691_),
    .B2(_08692_),
    .X(_08693_));
 sky130_fd_sc_hd__a2bb2o_2 _23024_ (.A1_N(_08688_),
    .A2_N(_08693_),
    .B1(_08688_),
    .B2(_08693_),
    .X(_08694_));
 sky130_fd_sc_hd__a2bb2o_2 _23025_ (.A1_N(_08687_),
    .A2_N(_08694_),
    .B1(_08687_),
    .B2(_08694_),
    .X(_08695_));
 sky130_fd_sc_hd__o22a_2 _23026_ (.A1(_08584_),
    .A2(_05169_),
    .B1(_06833_),
    .B2(_05845_),
    .X(_08696_));
 sky130_fd_sc_hd__and4_2 _23027_ (.A(_07680_),
    .B(_11923_),
    .C(_07681_),
    .D(_11920_),
    .X(_08697_));
 sky130_fd_sc_hd__nor2_2 _23028_ (.A(_08696_),
    .B(_08697_),
    .Y(_08698_));
 sky130_fd_sc_hd__nor2_2 _23029_ (.A(_07822_),
    .B(_05421_),
    .Y(_08699_));
 sky130_fd_sc_hd__a2bb2o_2 _23030_ (.A1_N(_08698_),
    .A2_N(_08699_),
    .B1(_08698_),
    .B2(_08699_),
    .X(_08700_));
 sky130_fd_sc_hd__or2_2 _23031_ (.A(_08098_),
    .B(_05937_),
    .X(_08701_));
 sky130_fd_sc_hd__and4_2 _23032_ (.A(_07686_),
    .B(_05014_),
    .C(_08100_),
    .D(_11926_),
    .X(_08702_));
 sky130_fd_sc_hd__o22a_2 _23033_ (.A1(_08592_),
    .A2(_11928_),
    .B1(_07545_),
    .B2(_05071_),
    .X(_08703_));
 sky130_fd_sc_hd__or2_2 _23034_ (.A(_08702_),
    .B(_08703_),
    .X(_08704_));
 sky130_fd_sc_hd__a2bb2o_2 _23035_ (.A1_N(_08701_),
    .A2_N(_08704_),
    .B1(_08701_),
    .B2(_08704_),
    .X(_08705_));
 sky130_fd_sc_hd__o21ba_2 _23036_ (.A1(_08590_),
    .A2(_08594_),
    .B1_N(_08591_),
    .X(_08706_));
 sky130_fd_sc_hd__a2bb2o_2 _23037_ (.A1_N(_08705_),
    .A2_N(_08706_),
    .B1(_08705_),
    .B2(_08706_),
    .X(_08707_));
 sky130_fd_sc_hd__a2bb2o_2 _23038_ (.A1_N(_08700_),
    .A2_N(_08707_),
    .B1(_08700_),
    .B2(_08707_),
    .X(_08708_));
 sky130_fd_sc_hd__o22a_2 _23039_ (.A1(_08595_),
    .A2(_08596_),
    .B1(_08589_),
    .B2(_08597_),
    .X(_08709_));
 sky130_fd_sc_hd__a2bb2o_2 _23040_ (.A1_N(_08708_),
    .A2_N(_08709_),
    .B1(_08708_),
    .B2(_08709_),
    .X(_08710_));
 sky130_fd_sc_hd__a2bb2o_2 _23041_ (.A1_N(_08695_),
    .A2_N(_08710_),
    .B1(_08695_),
    .B2(_08710_),
    .X(_08711_));
 sky130_fd_sc_hd__o22a_2 _23042_ (.A1(_08598_),
    .A2(_08599_),
    .B1(_08583_),
    .B2(_08600_),
    .X(_08712_));
 sky130_fd_sc_hd__a2bb2o_2 _23043_ (.A1_N(_08711_),
    .A2_N(_08712_),
    .B1(_08711_),
    .B2(_08712_),
    .X(_08713_));
 sky130_fd_sc_hd__a2bb2o_2 _23044_ (.A1_N(_08686_),
    .A2_N(_08713_),
    .B1(_08686_),
    .B2(_08713_),
    .X(_08714_));
 sky130_fd_sc_hd__o22a_2 _23045_ (.A1(_08601_),
    .A2(_08602_),
    .B1(_08574_),
    .B2(_08603_),
    .X(_08715_));
 sky130_fd_sc_hd__a2bb2o_2 _23046_ (.A1_N(_08714_),
    .A2_N(_08715_),
    .B1(_08714_),
    .B2(_08715_),
    .X(_08716_));
 sky130_fd_sc_hd__a2bb2o_2 _23047_ (.A1_N(_08669_),
    .A2_N(_08716_),
    .B1(_08669_),
    .B2(_08716_),
    .X(_08717_));
 sky130_fd_sc_hd__o22a_2 _23048_ (.A1(_08604_),
    .A2(_08605_),
    .B1(_08556_),
    .B2(_08606_),
    .X(_08718_));
 sky130_fd_sc_hd__a2bb2o_2 _23049_ (.A1_N(_08717_),
    .A2_N(_08718_),
    .B1(_08717_),
    .B2(_08718_),
    .X(_08719_));
 sky130_fd_sc_hd__a2bb2o_2 _23050_ (.A1_N(_08640_),
    .A2_N(_08719_),
    .B1(_08640_),
    .B2(_08719_),
    .X(_08720_));
 sky130_fd_sc_hd__o22a_2 _23051_ (.A1(_08607_),
    .A2(_08608_),
    .B1(_08525_),
    .B2(_08609_),
    .X(_08721_));
 sky130_fd_sc_hd__a2bb2o_2 _23052_ (.A1_N(_08720_),
    .A2_N(_08721_),
    .B1(_08720_),
    .B2(_08721_),
    .X(_08722_));
 sky130_fd_sc_hd__a2bb2o_2 _23053_ (.A1_N(_08622_),
    .A2_N(_08722_),
    .B1(_08622_),
    .B2(_08722_),
    .X(_08723_));
 sky130_fd_sc_hd__o22a_2 _23054_ (.A1(_08610_),
    .A2(_08611_),
    .B1(_08509_),
    .B2(_08612_),
    .X(_08724_));
 sky130_fd_sc_hd__a2bb2o_2 _23055_ (.A1_N(_08723_),
    .A2_N(_08724_),
    .B1(_08723_),
    .B2(_08724_),
    .X(_08725_));
 sky130_fd_sc_hd__a2bb2o_2 _23056_ (.A1_N(_08508_),
    .A2_N(_08725_),
    .B1(_08508_),
    .B2(_08725_),
    .X(_08726_));
 sky130_fd_sc_hd__o22a_2 _23057_ (.A1(_08613_),
    .A2(_08614_),
    .B1(_08376_),
    .B2(_08615_),
    .X(_08727_));
 sky130_fd_sc_hd__or2_2 _23058_ (.A(_08726_),
    .B(_08727_),
    .X(_08728_));
 sky130_fd_sc_hd__a21bo_2 _23059_ (.A1(_08726_),
    .A2(_08727_),
    .B1_N(_08728_),
    .X(_08729_));
 sky130_fd_sc_hd__a22o_2 _23060_ (.A1(_08506_),
    .A2(_08616_),
    .B1(_08495_),
    .B2(_08617_),
    .X(_08730_));
 sky130_fd_sc_hd__o31a_2 _23061_ (.A1(_08496_),
    .A2(_08618_),
    .A3(_08504_),
    .B1(_08730_),
    .X(_08731_));
 sky130_fd_sc_hd__a2bb2oi_2 _23062_ (.A1_N(_08729_),
    .A2_N(_08731_),
    .B1(_08729_),
    .B2(_08731_),
    .Y(_02661_));
 sky130_fd_sc_hd__o22a_2 _23063_ (.A1(_08723_),
    .A2(_08724_),
    .B1(_08508_),
    .B2(_08725_),
    .X(_08732_));
 sky130_fd_sc_hd__o22a_2 _23064_ (.A1(_08625_),
    .A2(_08638_),
    .B1(_08624_),
    .B2(_08639_),
    .X(_08733_));
 sky130_fd_sc_hd__or2_2 _23065_ (.A(_08373_),
    .B(_08733_),
    .X(_08734_));
 sky130_fd_sc_hd__a21bo_2 _23066_ (.A1(_08375_),
    .A2(_08733_),
    .B1_N(_08734_),
    .X(_08735_));
 sky130_fd_sc_hd__o22a_2 _23067_ (.A1(_08634_),
    .A2(_08635_),
    .B1(_08379_),
    .B2(_08637_),
    .X(_08736_));
 sky130_fd_sc_hd__o22a_2 _23068_ (.A1(_08642_),
    .A2(_08667_),
    .B1(_08641_),
    .B2(_08668_),
    .X(_08737_));
 sky130_fd_sc_hd__o22a_2 _23069_ (.A1(_08652_),
    .A2(_08653_),
    .B1(_08647_),
    .B2(_08654_),
    .X(_08738_));
 sky130_fd_sc_hd__o32a_2 _23070_ (.A1(_08038_),
    .A2(_08266_),
    .A3(_08644_),
    .B1(_08533_),
    .B2(_08646_),
    .X(_08739_));
 sky130_fd_sc_hd__a2bb2o_2 _23071_ (.A1_N(_08390_),
    .A2_N(_08739_),
    .B1(_08390_),
    .B2(_08739_),
    .X(_08740_));
 sky130_fd_sc_hd__a2bb2o_2 _23072_ (.A1_N(_08627_),
    .A2_N(_08740_),
    .B1(_08627_),
    .B2(_08740_),
    .X(_08741_));
 sky130_fd_sc_hd__o2bb2ai_2 _23073_ (.A1_N(_08738_),
    .A2_N(_08741_),
    .B1(_08738_),
    .B2(_08741_),
    .Y(_08742_));
 sky130_fd_sc_hd__buf_1 _23074_ (.A(_08627_),
    .X(_08743_));
 sky130_fd_sc_hd__o22a_2 _23075_ (.A1(_08389_),
    .A2(_08628_),
    .B1(_08743_),
    .B2(_08629_),
    .X(_08744_));
 sky130_fd_sc_hd__o2bb2a_2 _23076_ (.A1_N(_08742_),
    .A2_N(_08744_),
    .B1(_08742_),
    .B2(_08744_),
    .X(_08745_));
 sky130_vsdinv _23077_ (.A(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__o22a_2 _23078_ (.A1(_08626_),
    .A2(_08630_),
    .B1(_08631_),
    .B2(_08632_),
    .X(_08747_));
 sky130_vsdinv _23079_ (.A(_08747_),
    .Y(_08748_));
 sky130_fd_sc_hd__a22o_2 _23080_ (.A1(_08746_),
    .A2(_08747_),
    .B1(_08745_),
    .B2(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__a2bb2o_2 _23081_ (.A1_N(_08261_),
    .A2_N(_08749_),
    .B1(_08261_),
    .B2(_08749_),
    .X(_08750_));
 sky130_fd_sc_hd__a2bb2o_2 _23082_ (.A1_N(_08737_),
    .A2_N(_08750_),
    .B1(_08737_),
    .B2(_08750_),
    .X(_08751_));
 sky130_fd_sc_hd__a2bb2o_2 _23083_ (.A1_N(_08736_),
    .A2_N(_08751_),
    .B1(_08736_),
    .B2(_08751_),
    .X(_08752_));
 sky130_fd_sc_hd__o22a_2 _23084_ (.A1(_08664_),
    .A2(_08665_),
    .B1(_08655_),
    .B2(_08666_),
    .X(_08753_));
 sky130_fd_sc_hd__o22a_2 _23085_ (.A1(_08671_),
    .A2(_08684_),
    .B1(_08670_),
    .B2(_08685_),
    .X(_08754_));
 sky130_fd_sc_hd__or2_2 _23086_ (.A(_10584_),
    .B(_05007_),
    .X(_08755_));
 sky130_fd_sc_hd__a32o_2 _23087_ (.A1(_07868_),
    .A2(_05143_),
    .A3(_08645_),
    .B1(_08644_),
    .B2(_08755_),
    .X(_08756_));
 sky130_fd_sc_hd__a2bb2o_2 _23088_ (.A1_N(_08533_),
    .A2_N(_08756_),
    .B1(_08533_),
    .B2(_08756_),
    .X(_08757_));
 sky130_fd_sc_hd__buf_1 _23089_ (.A(_08757_),
    .X(_08758_));
 sky130_fd_sc_hd__o22a_2 _23090_ (.A1(_05405_),
    .A2(_06889_),
    .B1(_05131_),
    .B2(_07021_),
    .X(_08759_));
 sky130_fd_sc_hd__and4_2 _23091_ (.A(_11607_),
    .B(\pcpi_mul.rs1[29] ),
    .C(_11610_),
    .D(\pcpi_mul.rs1[30] ),
    .X(_08760_));
 sky130_fd_sc_hd__nor2_2 _23092_ (.A(_08759_),
    .B(_08760_),
    .Y(_08761_));
 sky130_fd_sc_hd__nor2_2 _23093_ (.A(_05057_),
    .B(_08266_),
    .Y(_08762_));
 sky130_fd_sc_hd__a2bb2o_2 _23094_ (.A1_N(_08761_),
    .A2_N(_08762_),
    .B1(_08761_),
    .B2(_08762_),
    .X(_08763_));
 sky130_fd_sc_hd__a21oi_2 _23095_ (.A1(_08650_),
    .A2(_08651_),
    .B1(_08649_),
    .Y(_08764_));
 sky130_fd_sc_hd__a2bb2o_2 _23096_ (.A1_N(_08763_),
    .A2_N(_08764_),
    .B1(_08763_),
    .B2(_08764_),
    .X(_08765_));
 sky130_fd_sc_hd__a2bb2o_2 _23097_ (.A1_N(_08758_),
    .A2_N(_08765_),
    .B1(_08758_),
    .B2(_08765_),
    .X(_08766_));
 sky130_fd_sc_hd__a21oi_2 _23098_ (.A1(_08660_),
    .A2(_08661_),
    .B1(_08659_),
    .Y(_08767_));
 sky130_fd_sc_hd__a21oi_2 _23099_ (.A1(_08674_),
    .A2(_08675_),
    .B1(_08673_),
    .Y(_08768_));
 sky130_fd_sc_hd__o22a_2 _23100_ (.A1(_08298_),
    .A2(_06742_),
    .B1(_08176_),
    .B2(_06878_),
    .X(_08769_));
 sky130_fd_sc_hd__and4_2 _23101_ (.A(_08300_),
    .B(_07459_),
    .C(_08301_),
    .D(_11884_),
    .X(_08770_));
 sky130_fd_sc_hd__nor2_2 _23102_ (.A(_08769_),
    .B(_08770_),
    .Y(_08771_));
 sky130_fd_sc_hd__nor2_2 _23103_ (.A(_07922_),
    .B(_06750_),
    .Y(_08772_));
 sky130_fd_sc_hd__a2bb2o_2 _23104_ (.A1_N(_08771_),
    .A2_N(_08772_),
    .B1(_08771_),
    .B2(_08772_),
    .X(_08773_));
 sky130_fd_sc_hd__a2bb2o_2 _23105_ (.A1_N(_08768_),
    .A2_N(_08773_),
    .B1(_08768_),
    .B2(_08773_),
    .X(_08774_));
 sky130_fd_sc_hd__a2bb2o_2 _23106_ (.A1_N(_08767_),
    .A2_N(_08774_),
    .B1(_08767_),
    .B2(_08774_),
    .X(_08775_));
 sky130_fd_sc_hd__o22a_2 _23107_ (.A1(_08657_),
    .A2(_08662_),
    .B1(_08656_),
    .B2(_08663_),
    .X(_08776_));
 sky130_fd_sc_hd__a2bb2o_2 _23108_ (.A1_N(_08775_),
    .A2_N(_08776_),
    .B1(_08775_),
    .B2(_08776_),
    .X(_08777_));
 sky130_fd_sc_hd__a2bb2o_2 _23109_ (.A1_N(_08766_),
    .A2_N(_08777_),
    .B1(_08766_),
    .B2(_08777_),
    .X(_08778_));
 sky130_fd_sc_hd__a2bb2o_2 _23110_ (.A1_N(_08754_),
    .A2_N(_08778_),
    .B1(_08754_),
    .B2(_08778_),
    .X(_08779_));
 sky130_fd_sc_hd__a2bb2o_2 _23111_ (.A1_N(_08753_),
    .A2_N(_08779_),
    .B1(_08753_),
    .B2(_08779_),
    .X(_08780_));
 sky130_fd_sc_hd__o22a_2 _23112_ (.A1(_08681_),
    .A2(_08682_),
    .B1(_08676_),
    .B2(_08683_),
    .X(_08781_));
 sky130_fd_sc_hd__o22a_2 _23113_ (.A1(_08688_),
    .A2(_08693_),
    .B1(_08687_),
    .B2(_08694_),
    .X(_08782_));
 sky130_fd_sc_hd__o22a_2 _23114_ (.A1(_07651_),
    .A2(_06359_),
    .B1(_08431_),
    .B2(_06361_),
    .X(_08783_));
 sky130_fd_sc_hd__and4_2 _23115_ (.A(_08433_),
    .B(_11897_),
    .C(_08434_),
    .D(_11895_),
    .X(_08784_));
 sky130_fd_sc_hd__nor2_2 _23116_ (.A(_08783_),
    .B(_08784_),
    .Y(_08785_));
 sky130_fd_sc_hd__nor2_2 _23117_ (.A(_08437_),
    .B(_06378_),
    .Y(_08786_));
 sky130_fd_sc_hd__a2bb2o_2 _23118_ (.A1_N(_08785_),
    .A2_N(_08786_),
    .B1(_08785_),
    .B2(_08786_),
    .X(_08787_));
 sky130_fd_sc_hd__o22a_2 _23119_ (.A1(_08440_),
    .A2(_05823_),
    .B1(_08441_),
    .B2(_06501_),
    .X(_08788_));
 sky130_fd_sc_hd__and4_2 _23120_ (.A(_07801_),
    .B(_11905_),
    .C(_07802_),
    .D(_11902_),
    .X(_08789_));
 sky130_fd_sc_hd__nor2_2 _23121_ (.A(_08788_),
    .B(_08789_),
    .Y(_08790_));
 sky130_fd_sc_hd__nor2_2 _23122_ (.A(_08445_),
    .B(_05996_),
    .Y(_08791_));
 sky130_fd_sc_hd__a2bb2o_2 _23123_ (.A1_N(_08790_),
    .A2_N(_08791_),
    .B1(_08790_),
    .B2(_08791_),
    .X(_08792_));
 sky130_fd_sc_hd__a21oi_2 _23124_ (.A1(_08679_),
    .A2(_08680_),
    .B1(_08678_),
    .Y(_08793_));
 sky130_fd_sc_hd__a2bb2o_2 _23125_ (.A1_N(_08792_),
    .A2_N(_08793_),
    .B1(_08792_),
    .B2(_08793_),
    .X(_08794_));
 sky130_fd_sc_hd__a2bb2o_2 _23126_ (.A1_N(_08787_),
    .A2_N(_08794_),
    .B1(_08787_),
    .B2(_08794_),
    .X(_08795_));
 sky130_fd_sc_hd__a2bb2o_2 _23127_ (.A1_N(_08782_),
    .A2_N(_08795_),
    .B1(_08782_),
    .B2(_08795_),
    .X(_08796_));
 sky130_fd_sc_hd__a2bb2o_2 _23128_ (.A1_N(_08781_),
    .A2_N(_08796_),
    .B1(_08781_),
    .B2(_08796_),
    .X(_08797_));
 sky130_fd_sc_hd__a21oi_2 _23129_ (.A1(_08691_),
    .A2(_08692_),
    .B1(_08690_),
    .Y(_08798_));
 sky130_fd_sc_hd__a21oi_2 _23130_ (.A1(_08698_),
    .A2(_08699_),
    .B1(_08697_),
    .Y(_08799_));
 sky130_fd_sc_hd__o22a_2 _23131_ (.A1(_07814_),
    .A2(_05598_),
    .B1(_06445_),
    .B2(_07059_),
    .X(_08800_));
 sky130_fd_sc_hd__and4_2 _23132_ (.A(_07816_),
    .B(_05897_),
    .C(_07672_),
    .D(_05999_),
    .X(_08801_));
 sky130_fd_sc_hd__nor2_2 _23133_ (.A(_08800_),
    .B(_08801_),
    .Y(_08802_));
 sky130_fd_sc_hd__nor2_2 _23134_ (.A(_06447_),
    .B(_05716_),
    .Y(_08803_));
 sky130_fd_sc_hd__a2bb2o_2 _23135_ (.A1_N(_08802_),
    .A2_N(_08803_),
    .B1(_08802_),
    .B2(_08803_),
    .X(_08804_));
 sky130_fd_sc_hd__a2bb2o_2 _23136_ (.A1_N(_08799_),
    .A2_N(_08804_),
    .B1(_08799_),
    .B2(_08804_),
    .X(_08805_));
 sky130_fd_sc_hd__a2bb2o_2 _23137_ (.A1_N(_08798_),
    .A2_N(_08805_),
    .B1(_08798_),
    .B2(_08805_),
    .X(_08806_));
 sky130_fd_sc_hd__o22a_2 _23138_ (.A1(_08584_),
    .A2(_05256_),
    .B1(_06833_),
    .B2(_05720_),
    .X(_08807_));
 sky130_fd_sc_hd__and4_2 _23139_ (.A(_07680_),
    .B(_11920_),
    .C(_07681_),
    .D(_11917_),
    .X(_08808_));
 sky130_fd_sc_hd__nor2_2 _23140_ (.A(_08807_),
    .B(_08808_),
    .Y(_08809_));
 sky130_fd_sc_hd__nor2_2 _23141_ (.A(_07822_),
    .B(_05502_),
    .Y(_08810_));
 sky130_fd_sc_hd__a2bb2o_2 _23142_ (.A1_N(_08809_),
    .A2_N(_08810_),
    .B1(_08809_),
    .B2(_08810_),
    .X(_08811_));
 sky130_fd_sc_hd__or2_2 _23143_ (.A(_08098_),
    .B(_05169_),
    .X(_08812_));
 sky130_fd_sc_hd__and4_2 _23144_ (.A(_07686_),
    .B(_05071_),
    .C(_11559_),
    .D(_11924_),
    .X(_08813_));
 sky130_fd_sc_hd__o22a_2 _23145_ (.A1(_08592_),
    .A2(_11926_),
    .B1(_07545_),
    .B2(_05081_),
    .X(_08814_));
 sky130_fd_sc_hd__or2_2 _23146_ (.A(_08813_),
    .B(_08814_),
    .X(_08815_));
 sky130_fd_sc_hd__a2bb2o_2 _23147_ (.A1_N(_08812_),
    .A2_N(_08815_),
    .B1(_08812_),
    .B2(_08815_),
    .X(_08816_));
 sky130_fd_sc_hd__o21ba_2 _23148_ (.A1(_08701_),
    .A2(_08704_),
    .B1_N(_08702_),
    .X(_08817_));
 sky130_fd_sc_hd__a2bb2o_2 _23149_ (.A1_N(_08816_),
    .A2_N(_08817_),
    .B1(_08816_),
    .B2(_08817_),
    .X(_08818_));
 sky130_fd_sc_hd__a2bb2o_2 _23150_ (.A1_N(_08811_),
    .A2_N(_08818_),
    .B1(_08811_),
    .B2(_08818_),
    .X(_08819_));
 sky130_fd_sc_hd__o22a_2 _23151_ (.A1(_08705_),
    .A2(_08706_),
    .B1(_08700_),
    .B2(_08707_),
    .X(_08820_));
 sky130_fd_sc_hd__a2bb2o_2 _23152_ (.A1_N(_08819_),
    .A2_N(_08820_),
    .B1(_08819_),
    .B2(_08820_),
    .X(_08821_));
 sky130_fd_sc_hd__a2bb2o_2 _23153_ (.A1_N(_08806_),
    .A2_N(_08821_),
    .B1(_08806_),
    .B2(_08821_),
    .X(_08822_));
 sky130_fd_sc_hd__o22a_2 _23154_ (.A1(_08708_),
    .A2(_08709_),
    .B1(_08695_),
    .B2(_08710_),
    .X(_08823_));
 sky130_fd_sc_hd__a2bb2o_2 _23155_ (.A1_N(_08822_),
    .A2_N(_08823_),
    .B1(_08822_),
    .B2(_08823_),
    .X(_08824_));
 sky130_fd_sc_hd__a2bb2o_2 _23156_ (.A1_N(_08797_),
    .A2_N(_08824_),
    .B1(_08797_),
    .B2(_08824_),
    .X(_08825_));
 sky130_fd_sc_hd__o22a_2 _23157_ (.A1(_08711_),
    .A2(_08712_),
    .B1(_08686_),
    .B2(_08713_),
    .X(_08826_));
 sky130_fd_sc_hd__a2bb2o_2 _23158_ (.A1_N(_08825_),
    .A2_N(_08826_),
    .B1(_08825_),
    .B2(_08826_),
    .X(_08827_));
 sky130_fd_sc_hd__a2bb2o_2 _23159_ (.A1_N(_08780_),
    .A2_N(_08827_),
    .B1(_08780_),
    .B2(_08827_),
    .X(_08828_));
 sky130_fd_sc_hd__o22a_2 _23160_ (.A1(_08714_),
    .A2(_08715_),
    .B1(_08669_),
    .B2(_08716_),
    .X(_08829_));
 sky130_fd_sc_hd__a2bb2o_2 _23161_ (.A1_N(_08828_),
    .A2_N(_08829_),
    .B1(_08828_),
    .B2(_08829_),
    .X(_08830_));
 sky130_fd_sc_hd__a2bb2o_2 _23162_ (.A1_N(_08752_),
    .A2_N(_08830_),
    .B1(_08752_),
    .B2(_08830_),
    .X(_08831_));
 sky130_fd_sc_hd__o22a_2 _23163_ (.A1(_08717_),
    .A2(_08718_),
    .B1(_08640_),
    .B2(_08719_),
    .X(_08832_));
 sky130_fd_sc_hd__a2bb2o_2 _23164_ (.A1_N(_08831_),
    .A2_N(_08832_),
    .B1(_08831_),
    .B2(_08832_),
    .X(_08833_));
 sky130_fd_sc_hd__a2bb2o_2 _23165_ (.A1_N(_08735_),
    .A2_N(_08833_),
    .B1(_08735_),
    .B2(_08833_),
    .X(_08834_));
 sky130_fd_sc_hd__o22a_2 _23166_ (.A1(_08720_),
    .A2(_08721_),
    .B1(_08622_),
    .B2(_08722_),
    .X(_08835_));
 sky130_fd_sc_hd__a2bb2o_2 _23167_ (.A1_N(_08834_),
    .A2_N(_08835_),
    .B1(_08834_),
    .B2(_08835_),
    .X(_08836_));
 sky130_fd_sc_hd__a2bb2o_2 _23168_ (.A1_N(_08621_),
    .A2_N(_08836_),
    .B1(_08621_),
    .B2(_08836_),
    .X(_08837_));
 sky130_fd_sc_hd__and2_2 _23169_ (.A(_08732_),
    .B(_08837_),
    .X(_08838_));
 sky130_fd_sc_hd__or2_2 _23170_ (.A(_08732_),
    .B(_08837_),
    .X(_08839_));
 sky130_fd_sc_hd__or2b_2 _23171_ (.A(_08838_),
    .B_N(_08839_),
    .X(_08840_));
 sky130_fd_sc_hd__o21ai_2 _23172_ (.A1(_08729_),
    .A2(_08731_),
    .B1(_08728_),
    .Y(_08841_));
 sky130_fd_sc_hd__a2bb2o_2 _23173_ (.A1_N(_08840_),
    .A2_N(_08841_),
    .B1(_08840_),
    .B2(_08841_),
    .X(_02662_));
 sky130_fd_sc_hd__buf_1 _23174_ (.A(_08374_),
    .X(_08842_));
 sky130_fd_sc_hd__o22a_2 _23175_ (.A1(_08737_),
    .A2(_08750_),
    .B1(_08736_),
    .B2(_08751_),
    .X(_08843_));
 sky130_fd_sc_hd__or2_2 _23176_ (.A(_08374_),
    .B(_08843_),
    .X(_08844_));
 sky130_fd_sc_hd__a21bo_2 _23177_ (.A1(_08842_),
    .A2(_08843_),
    .B1_N(_08844_),
    .X(_08845_));
 sky130_fd_sc_hd__o22a_2 _23178_ (.A1(_08746_),
    .A2(_08747_),
    .B1(_08379_),
    .B2(_08749_),
    .X(_08846_));
 sky130_fd_sc_hd__o22a_2 _23179_ (.A1(_08754_),
    .A2(_08778_),
    .B1(_08753_),
    .B2(_08779_),
    .X(_08847_));
 sky130_fd_sc_hd__o22a_2 _23180_ (.A1(_08763_),
    .A2(_08764_),
    .B1(_08757_),
    .B2(_08765_),
    .X(_08848_));
 sky130_fd_sc_hd__o22a_2 _23181_ (.A1(_08644_),
    .A2(_08755_),
    .B1(_08532_),
    .B2(_08756_),
    .X(_08849_));
 sky130_fd_sc_hd__or2_2 _23182_ (.A(_08388_),
    .B(_08849_),
    .X(_08850_));
 sky130_fd_sc_hd__a21bo_2 _23183_ (.A1(_08388_),
    .A2(_08849_),
    .B1_N(_08850_),
    .X(_08851_));
 sky130_fd_sc_hd__a2bb2o_2 _23184_ (.A1_N(_08515_),
    .A2_N(_08851_),
    .B1(_08515_),
    .B2(_08851_),
    .X(_08852_));
 sky130_fd_sc_hd__buf_1 _23185_ (.A(_08852_),
    .X(_08853_));
 sky130_fd_sc_hd__o2bb2ai_2 _23186_ (.A1_N(_08848_),
    .A2_N(_08853_),
    .B1(_08848_),
    .B2(_08852_),
    .Y(_08854_));
 sky130_fd_sc_hd__o22a_2 _23187_ (.A1(_08389_),
    .A2(_08739_),
    .B1(_08743_),
    .B2(_08740_),
    .X(_08855_));
 sky130_fd_sc_hd__o2bb2a_2 _23188_ (.A1_N(_08854_),
    .A2_N(_08855_),
    .B1(_08854_),
    .B2(_08855_),
    .X(_08856_));
 sky130_vsdinv _23189_ (.A(_08856_),
    .Y(_08857_));
 sky130_fd_sc_hd__o22a_2 _23190_ (.A1(_08738_),
    .A2(_08741_),
    .B1(_08742_),
    .B2(_08744_),
    .X(_08858_));
 sky130_vsdinv _23191_ (.A(_08858_),
    .Y(_08859_));
 sky130_fd_sc_hd__a22o_2 _23192_ (.A1(_08857_),
    .A2(_08858_),
    .B1(_08856_),
    .B2(_08859_),
    .X(_08860_));
 sky130_fd_sc_hd__a2bb2o_2 _23193_ (.A1_N(_08512_),
    .A2_N(_08860_),
    .B1(_08512_),
    .B2(_08860_),
    .X(_08861_));
 sky130_fd_sc_hd__a2bb2o_2 _23194_ (.A1_N(_08847_),
    .A2_N(_08861_),
    .B1(_08847_),
    .B2(_08861_),
    .X(_08862_));
 sky130_fd_sc_hd__a2bb2o_2 _23195_ (.A1_N(_08846_),
    .A2_N(_08862_),
    .B1(_08846_),
    .B2(_08862_),
    .X(_08863_));
 sky130_fd_sc_hd__o22a_2 _23196_ (.A1(_08775_),
    .A2(_08776_),
    .B1(_08766_),
    .B2(_08777_),
    .X(_08864_));
 sky130_fd_sc_hd__o22a_2 _23197_ (.A1(_08782_),
    .A2(_08795_),
    .B1(_08781_),
    .B2(_08796_),
    .X(_08865_));
 sky130_fd_sc_hd__o22a_2 _23198_ (.A1(_05405_),
    .A2(_07021_),
    .B1(_05131_),
    .B2(_07732_),
    .X(_08866_));
 sky130_fd_sc_hd__and4_2 _23199_ (.A(_06928_),
    .B(\pcpi_mul.rs1[30] ),
    .C(_06929_),
    .D(\pcpi_mul.rs1[31] ),
    .X(_08867_));
 sky130_fd_sc_hd__nor2_2 _23200_ (.A(_08866_),
    .B(_08867_),
    .Y(_08868_));
 sky130_fd_sc_hd__nor2_2 _23201_ (.A(_07727_),
    .B(_05133_),
    .Y(_08869_));
 sky130_fd_sc_hd__a2bb2o_2 _23202_ (.A1_N(_08868_),
    .A2_N(_08869_),
    .B1(_08868_),
    .B2(_08869_),
    .X(_08870_));
 sky130_fd_sc_hd__a31o_2 _23203_ (.A1(\pcpi_mul.rs2[12] ),
    .A2(_11873_),
    .A3(_08761_),
    .B1(_08760_),
    .X(_08871_));
 sky130_vsdinv _23204_ (.A(_08871_),
    .Y(_08872_));
 sky130_vsdinv _23205_ (.A(_08870_),
    .Y(_08873_));
 sky130_fd_sc_hd__a22o_2 _23206_ (.A1(_08870_),
    .A2(_08872_),
    .B1(_08873_),
    .B2(_08871_),
    .X(_08874_));
 sky130_fd_sc_hd__a2bb2o_2 _23207_ (.A1_N(_08758_),
    .A2_N(_08874_),
    .B1(_08758_),
    .B2(_08874_),
    .X(_08875_));
 sky130_fd_sc_hd__a21oi_2 _23208_ (.A1(_08771_),
    .A2(_08772_),
    .B1(_08770_),
    .Y(_08876_));
 sky130_fd_sc_hd__a21oi_2 _23209_ (.A1(_08785_),
    .A2(_08786_),
    .B1(_08784_),
    .Y(_08877_));
 sky130_fd_sc_hd__o22a_2 _23210_ (.A1(_08298_),
    .A2(_06878_),
    .B1(_08176_),
    .B2(_06749_),
    .X(_08878_));
 sky130_fd_sc_hd__and4_2 _23211_ (.A(_08300_),
    .B(_11884_),
    .C(_08301_),
    .D(_07749_),
    .X(_08879_));
 sky130_fd_sc_hd__nor2_2 _23212_ (.A(_08878_),
    .B(_08879_),
    .Y(_08880_));
 sky130_fd_sc_hd__nor2_2 _23213_ (.A(_07346_),
    .B(_06891_),
    .Y(_08881_));
 sky130_fd_sc_hd__a2bb2o_2 _23214_ (.A1_N(_08880_),
    .A2_N(_08881_),
    .B1(_08880_),
    .B2(_08881_),
    .X(_08882_));
 sky130_fd_sc_hd__a2bb2o_2 _23215_ (.A1_N(_08877_),
    .A2_N(_08882_),
    .B1(_08877_),
    .B2(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__a2bb2o_2 _23216_ (.A1_N(_08876_),
    .A2_N(_08883_),
    .B1(_08876_),
    .B2(_08883_),
    .X(_08884_));
 sky130_fd_sc_hd__o22a_2 _23217_ (.A1(_08768_),
    .A2(_08773_),
    .B1(_08767_),
    .B2(_08774_),
    .X(_08885_));
 sky130_fd_sc_hd__a2bb2o_2 _23218_ (.A1_N(_08884_),
    .A2_N(_08885_),
    .B1(_08884_),
    .B2(_08885_),
    .X(_08886_));
 sky130_fd_sc_hd__a2bb2o_2 _23219_ (.A1_N(_08875_),
    .A2_N(_08886_),
    .B1(_08875_),
    .B2(_08886_),
    .X(_08887_));
 sky130_fd_sc_hd__a2bb2o_2 _23220_ (.A1_N(_08865_),
    .A2_N(_08887_),
    .B1(_08865_),
    .B2(_08887_),
    .X(_08888_));
 sky130_fd_sc_hd__a2bb2o_2 _23221_ (.A1_N(_08864_),
    .A2_N(_08888_),
    .B1(_08864_),
    .B2(_08888_),
    .X(_08889_));
 sky130_fd_sc_hd__o22a_2 _23222_ (.A1(_08792_),
    .A2(_08793_),
    .B1(_08787_),
    .B2(_08794_),
    .X(_08890_));
 sky130_fd_sc_hd__o22a_2 _23223_ (.A1(_08799_),
    .A2(_08804_),
    .B1(_08798_),
    .B2(_08805_),
    .X(_08891_));
 sky130_fd_sc_hd__o22a_2 _23224_ (.A1(_07651_),
    .A2(_06361_),
    .B1(_05659_),
    .B2(_06616_),
    .X(_08892_));
 sky130_fd_sc_hd__and4_2 _23225_ (.A(_11593_),
    .B(_11895_),
    .C(_08434_),
    .D(_06885_),
    .X(_08893_));
 sky130_fd_sc_hd__nor2_2 _23226_ (.A(_08892_),
    .B(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__nor2_2 _23227_ (.A(_05562_),
    .B(_06497_),
    .Y(_08895_));
 sky130_fd_sc_hd__a2bb2o_2 _23228_ (.A1_N(_08894_),
    .A2_N(_08895_),
    .B1(_08894_),
    .B2(_08895_),
    .X(_08896_));
 sky130_fd_sc_hd__o22a_2 _23229_ (.A1(_08440_),
    .A2(_06501_),
    .B1(_06034_),
    .B2(_06904_),
    .X(_08897_));
 sky130_fd_sc_hd__and4_2 _23230_ (.A(_07801_),
    .B(_11902_),
    .C(_07802_),
    .D(_06499_),
    .X(_08898_));
 sky130_fd_sc_hd__nor2_2 _23231_ (.A(_08897_),
    .B(_08898_),
    .Y(_08899_));
 sky130_fd_sc_hd__nor2_2 _23232_ (.A(_08445_),
    .B(_06112_),
    .Y(_08900_));
 sky130_fd_sc_hd__a2bb2o_2 _23233_ (.A1_N(_08899_),
    .A2_N(_08900_),
    .B1(_08899_),
    .B2(_08900_),
    .X(_08901_));
 sky130_fd_sc_hd__a21oi_2 _23234_ (.A1(_08790_),
    .A2(_08791_),
    .B1(_08789_),
    .Y(_08902_));
 sky130_fd_sc_hd__a2bb2o_2 _23235_ (.A1_N(_08901_),
    .A2_N(_08902_),
    .B1(_08901_),
    .B2(_08902_),
    .X(_08903_));
 sky130_fd_sc_hd__a2bb2o_2 _23236_ (.A1_N(_08896_),
    .A2_N(_08903_),
    .B1(_08896_),
    .B2(_08903_),
    .X(_08904_));
 sky130_fd_sc_hd__a2bb2o_2 _23237_ (.A1_N(_08891_),
    .A2_N(_08904_),
    .B1(_08891_),
    .B2(_08904_),
    .X(_08905_));
 sky130_fd_sc_hd__a2bb2o_2 _23238_ (.A1_N(_08890_),
    .A2_N(_08905_),
    .B1(_08890_),
    .B2(_08905_),
    .X(_08906_));
 sky130_fd_sc_hd__a21oi_2 _23239_ (.A1(_08802_),
    .A2(_08803_),
    .B1(_08801_),
    .Y(_08907_));
 sky130_fd_sc_hd__a21oi_2 _23240_ (.A1(_08809_),
    .A2(_08810_),
    .B1(_08808_),
    .Y(_08908_));
 sky130_fd_sc_hd__buf_1 _23241_ (.A(_06974_),
    .X(_08909_));
 sky130_fd_sc_hd__o22a_2 _23242_ (.A1(_08909_),
    .A2(_07059_),
    .B1(_06442_),
    .B2(_07196_),
    .X(_08910_));
 sky130_fd_sc_hd__and4_2 _23243_ (.A(_11575_),
    .B(_05999_),
    .C(_08456_),
    .D(_06117_),
    .X(_08911_));
 sky130_fd_sc_hd__nor2_2 _23244_ (.A(_08910_),
    .B(_08911_),
    .Y(_08912_));
 sky130_fd_sc_hd__nor2_2 _23245_ (.A(_06273_),
    .B(_05885_),
    .Y(_08913_));
 sky130_fd_sc_hd__a2bb2o_2 _23246_ (.A1_N(_08912_),
    .A2_N(_08913_),
    .B1(_08912_),
    .B2(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__a2bb2o_2 _23247_ (.A1_N(_08908_),
    .A2_N(_08914_),
    .B1(_08908_),
    .B2(_08914_),
    .X(_08915_));
 sky130_fd_sc_hd__a2bb2o_2 _23248_ (.A1_N(_08907_),
    .A2_N(_08915_),
    .B1(_08907_),
    .B2(_08915_),
    .X(_08916_));
 sky130_fd_sc_hd__buf_1 _23249_ (.A(_07387_),
    .X(_08917_));
 sky130_fd_sc_hd__o22a_2 _23250_ (.A1(_08917_),
    .A2(_05343_),
    .B1(_06830_),
    .B2(_05828_),
    .X(_08918_));
 sky130_fd_sc_hd__and4_2 _23251_ (.A(_11567_),
    .B(_11917_),
    .C(_11571_),
    .D(_11915_),
    .X(_08919_));
 sky130_fd_sc_hd__nor2_2 _23252_ (.A(_08918_),
    .B(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__nor2_2 _23253_ (.A(_06687_),
    .B(_05599_),
    .Y(_08921_));
 sky130_fd_sc_hd__a2bb2o_2 _23254_ (.A1_N(_08920_),
    .A2_N(_08921_),
    .B1(_08920_),
    .B2(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__or2_2 _23255_ (.A(_08098_),
    .B(_05256_),
    .X(_08923_));
 sky130_fd_sc_hd__and4_2 _23256_ (.A(_07686_),
    .B(_05081_),
    .C(_08100_),
    .D(_11922_),
    .X(_08924_));
 sky130_fd_sc_hd__o22a_2 _23257_ (.A1(_08592_),
    .A2(_11924_),
    .B1(_07965_),
    .B2(_05168_),
    .X(_08925_));
 sky130_fd_sc_hd__or2_2 _23258_ (.A(_08924_),
    .B(_08925_),
    .X(_08926_));
 sky130_fd_sc_hd__a2bb2o_2 _23259_ (.A1_N(_08923_),
    .A2_N(_08926_),
    .B1(_08923_),
    .B2(_08926_),
    .X(_08927_));
 sky130_fd_sc_hd__o21ba_2 _23260_ (.A1(_08812_),
    .A2(_08815_),
    .B1_N(_08813_),
    .X(_08928_));
 sky130_fd_sc_hd__a2bb2o_2 _23261_ (.A1_N(_08927_),
    .A2_N(_08928_),
    .B1(_08927_),
    .B2(_08928_),
    .X(_08929_));
 sky130_fd_sc_hd__a2bb2o_2 _23262_ (.A1_N(_08922_),
    .A2_N(_08929_),
    .B1(_08922_),
    .B2(_08929_),
    .X(_08930_));
 sky130_fd_sc_hd__o22a_2 _23263_ (.A1(_08816_),
    .A2(_08817_),
    .B1(_08811_),
    .B2(_08818_),
    .X(_08931_));
 sky130_fd_sc_hd__a2bb2o_2 _23264_ (.A1_N(_08930_),
    .A2_N(_08931_),
    .B1(_08930_),
    .B2(_08931_),
    .X(_08932_));
 sky130_fd_sc_hd__a2bb2o_2 _23265_ (.A1_N(_08916_),
    .A2_N(_08932_),
    .B1(_08916_),
    .B2(_08932_),
    .X(_08933_));
 sky130_fd_sc_hd__o22a_2 _23266_ (.A1(_08819_),
    .A2(_08820_),
    .B1(_08806_),
    .B2(_08821_),
    .X(_08934_));
 sky130_fd_sc_hd__a2bb2o_2 _23267_ (.A1_N(_08933_),
    .A2_N(_08934_),
    .B1(_08933_),
    .B2(_08934_),
    .X(_08935_));
 sky130_fd_sc_hd__a2bb2o_2 _23268_ (.A1_N(_08906_),
    .A2_N(_08935_),
    .B1(_08906_),
    .B2(_08935_),
    .X(_08936_));
 sky130_fd_sc_hd__o22a_2 _23269_ (.A1(_08822_),
    .A2(_08823_),
    .B1(_08797_),
    .B2(_08824_),
    .X(_08937_));
 sky130_fd_sc_hd__a2bb2o_2 _23270_ (.A1_N(_08936_),
    .A2_N(_08937_),
    .B1(_08936_),
    .B2(_08937_),
    .X(_08938_));
 sky130_fd_sc_hd__a2bb2o_2 _23271_ (.A1_N(_08889_),
    .A2_N(_08938_),
    .B1(_08889_),
    .B2(_08938_),
    .X(_08939_));
 sky130_fd_sc_hd__o22a_2 _23272_ (.A1(_08825_),
    .A2(_08826_),
    .B1(_08780_),
    .B2(_08827_),
    .X(_08940_));
 sky130_fd_sc_hd__a2bb2o_2 _23273_ (.A1_N(_08939_),
    .A2_N(_08940_),
    .B1(_08939_),
    .B2(_08940_),
    .X(_08941_));
 sky130_fd_sc_hd__a2bb2o_2 _23274_ (.A1_N(_08863_),
    .A2_N(_08941_),
    .B1(_08863_),
    .B2(_08941_),
    .X(_08942_));
 sky130_fd_sc_hd__o22a_2 _23275_ (.A1(_08828_),
    .A2(_08829_),
    .B1(_08752_),
    .B2(_08830_),
    .X(_08943_));
 sky130_fd_sc_hd__a2bb2o_2 _23276_ (.A1_N(_08942_),
    .A2_N(_08943_),
    .B1(_08942_),
    .B2(_08943_),
    .X(_08944_));
 sky130_fd_sc_hd__a2bb2o_2 _23277_ (.A1_N(_08845_),
    .A2_N(_08944_),
    .B1(_08845_),
    .B2(_08944_),
    .X(_08945_));
 sky130_fd_sc_hd__o22a_2 _23278_ (.A1(_08831_),
    .A2(_08832_),
    .B1(_08735_),
    .B2(_08833_),
    .X(_08946_));
 sky130_fd_sc_hd__a2bb2o_2 _23279_ (.A1_N(_08945_),
    .A2_N(_08946_),
    .B1(_08945_),
    .B2(_08946_),
    .X(_08947_));
 sky130_fd_sc_hd__a2bb2o_2 _23280_ (.A1_N(_08734_),
    .A2_N(_08947_),
    .B1(_08734_),
    .B2(_08947_),
    .X(_08948_));
 sky130_fd_sc_hd__o22a_2 _23281_ (.A1(_08834_),
    .A2(_08835_),
    .B1(_08621_),
    .B2(_08836_),
    .X(_08949_));
 sky130_fd_sc_hd__or2_2 _23282_ (.A(_08948_),
    .B(_08949_),
    .X(_08950_));
 sky130_fd_sc_hd__a21bo_2 _23283_ (.A1(_08948_),
    .A2(_08949_),
    .B1_N(_08950_),
    .X(_08951_));
 sky130_fd_sc_hd__or2_2 _23284_ (.A(_08729_),
    .B(_08840_),
    .X(_08952_));
 sky130_fd_sc_hd__or3_2 _23285_ (.A(_08496_),
    .B(_08618_),
    .C(_08952_),
    .X(_08953_));
 sky130_fd_sc_hd__o221a_2 _23286_ (.A1(_08728_),
    .A2(_08838_),
    .B1(_08730_),
    .B2(_08952_),
    .C1(_08839_),
    .X(_08954_));
 sky130_fd_sc_hd__o21ai_2 _23287_ (.A1(_08504_),
    .A2(_08953_),
    .B1(_08954_),
    .Y(_08955_));
 sky130_vsdinv _23288_ (.A(_08955_),
    .Y(_08956_));
 sky130_vsdinv _23289_ (.A(_08951_),
    .Y(_08957_));
 sky130_fd_sc_hd__o22a_2 _23290_ (.A1(_08951_),
    .A2(_08956_),
    .B1(_08957_),
    .B2(_08955_),
    .X(_02663_));
 sky130_fd_sc_hd__o22a_2 _23291_ (.A1(_08945_),
    .A2(_08946_),
    .B1(_08734_),
    .B2(_08947_),
    .X(_08958_));
 sky130_fd_sc_hd__o22a_2 _23292_ (.A1(_08847_),
    .A2(_08861_),
    .B1(_08846_),
    .B2(_08862_),
    .X(_08959_));
 sky130_fd_sc_hd__or2_2 _23293_ (.A(_08373_),
    .B(_08959_),
    .X(_08960_));
 sky130_fd_sc_hd__a21bo_2 _23294_ (.A1(_08375_),
    .A2(_08959_),
    .B1_N(_08960_),
    .X(_08961_));
 sky130_fd_sc_hd__o22a_2 _23295_ (.A1(_08857_),
    .A2(_08858_),
    .B1(_08623_),
    .B2(_08860_),
    .X(_08962_));
 sky130_fd_sc_hd__o22a_2 _23296_ (.A1(_08865_),
    .A2(_08887_),
    .B1(_08864_),
    .B2(_08888_),
    .X(_08963_));
 sky130_fd_sc_hd__o22a_2 _23297_ (.A1(_08870_),
    .A2(_08872_),
    .B1(_08757_),
    .B2(_08874_),
    .X(_08964_));
 sky130_fd_sc_hd__a2bb2o_2 _23298_ (.A1_N(_08852_),
    .A2_N(_08964_),
    .B1(_08852_),
    .B2(_08964_),
    .X(_08965_));
 sky130_fd_sc_hd__o21a_2 _23299_ (.A1(_08743_),
    .A2(_08851_),
    .B1(_08850_),
    .X(_08966_));
 sky130_fd_sc_hd__o2bb2a_2 _23300_ (.A1_N(_08965_),
    .A2_N(_08966_),
    .B1(_08965_),
    .B2(_08966_),
    .X(_08967_));
 sky130_vsdinv _23301_ (.A(_08967_),
    .Y(_08968_));
 sky130_fd_sc_hd__o22a_2 _23302_ (.A1(_08848_),
    .A2(_08853_),
    .B1(_08854_),
    .B2(_08855_),
    .X(_08969_));
 sky130_vsdinv _23303_ (.A(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__a22o_2 _23304_ (.A1(_08968_),
    .A2(_08969_),
    .B1(_08967_),
    .B2(_08970_),
    .X(_08971_));
 sky130_fd_sc_hd__a2bb2o_2 _23305_ (.A1_N(_08512_),
    .A2_N(_08971_),
    .B1(_08512_),
    .B2(_08971_),
    .X(_08972_));
 sky130_fd_sc_hd__a2bb2o_2 _23306_ (.A1_N(_08963_),
    .A2_N(_08972_),
    .B1(_08963_),
    .B2(_08972_),
    .X(_08973_));
 sky130_fd_sc_hd__a2bb2o_2 _23307_ (.A1_N(_08962_),
    .A2_N(_08973_),
    .B1(_08962_),
    .B2(_08973_),
    .X(_08974_));
 sky130_fd_sc_hd__o22a_2 _23308_ (.A1(_08884_),
    .A2(_08885_),
    .B1(_08875_),
    .B2(_08886_),
    .X(_08975_));
 sky130_fd_sc_hd__o22a_2 _23309_ (.A1(_08891_),
    .A2(_08904_),
    .B1(_08890_),
    .B2(_08905_),
    .X(_08976_));
 sky130_fd_sc_hd__a31o_2 _23310_ (.A1(_07869_),
    .A2(\pcpi_mul.rs2[12] ),
    .A3(_08868_),
    .B1(_08867_),
    .X(_08977_));
 sky130_vsdinv _23311_ (.A(_08977_),
    .Y(_08978_));
 sky130_fd_sc_hd__o22a_2 _23312_ (.A1(_07626_),
    .A2(_07159_),
    .B1(_07727_),
    .B2(_05132_),
    .X(_08979_));
 sky130_fd_sc_hd__and4_2 _23313_ (.A(_11608_),
    .B(_11873_),
    .C(_07868_),
    .D(_11611_),
    .X(_08980_));
 sky130_fd_sc_hd__nor2_2 _23314_ (.A(_08979_),
    .B(_08980_),
    .Y(_08981_));
 sky130_fd_sc_hd__o2bb2a_2 _23315_ (.A1_N(_08869_),
    .A2_N(_08981_),
    .B1(_08869_),
    .B2(_08981_),
    .X(_08982_));
 sky130_vsdinv _23316_ (.A(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__a22o_2 _23317_ (.A1(_08978_),
    .A2(_08983_),
    .B1(_08977_),
    .B2(_08982_),
    .X(_08984_));
 sky130_fd_sc_hd__a2bb2o_2 _23318_ (.A1_N(_08758_),
    .A2_N(_08984_),
    .B1(_08758_),
    .B2(_08984_),
    .X(_08985_));
 sky130_fd_sc_hd__a21oi_2 _23319_ (.A1(_08880_),
    .A2(_08881_),
    .B1(_08879_),
    .Y(_08986_));
 sky130_fd_sc_hd__a21oi_2 _23320_ (.A1(_08894_),
    .A2(_08895_),
    .B1(_08893_),
    .Y(_08987_));
 sky130_fd_sc_hd__o22a_2 _23321_ (.A1(_07340_),
    .A2(_06749_),
    .B1(_05392_),
    .B2(_06890_),
    .X(_08988_));
 sky130_fd_sc_hd__and4_2 _23322_ (.A(_07342_),
    .B(_07749_),
    .C(_07343_),
    .D(_07587_),
    .X(_08989_));
 sky130_fd_sc_hd__nor2_2 _23323_ (.A(_08988_),
    .B(_08989_),
    .Y(_08990_));
 sky130_fd_sc_hd__nor2_2 _23324_ (.A(_07346_),
    .B(_07285_),
    .Y(_08991_));
 sky130_fd_sc_hd__a2bb2o_2 _23325_ (.A1_N(_08990_),
    .A2_N(_08991_),
    .B1(_08990_),
    .B2(_08991_),
    .X(_08992_));
 sky130_fd_sc_hd__a2bb2o_2 _23326_ (.A1_N(_08987_),
    .A2_N(_08992_),
    .B1(_08987_),
    .B2(_08992_),
    .X(_08993_));
 sky130_fd_sc_hd__a2bb2o_2 _23327_ (.A1_N(_08986_),
    .A2_N(_08993_),
    .B1(_08986_),
    .B2(_08993_),
    .X(_08994_));
 sky130_fd_sc_hd__o22a_2 _23328_ (.A1(_08877_),
    .A2(_08882_),
    .B1(_08876_),
    .B2(_08883_),
    .X(_08995_));
 sky130_fd_sc_hd__a2bb2o_2 _23329_ (.A1_N(_08994_),
    .A2_N(_08995_),
    .B1(_08994_),
    .B2(_08995_),
    .X(_08996_));
 sky130_fd_sc_hd__a2bb2o_2 _23330_ (.A1_N(_08985_),
    .A2_N(_08996_),
    .B1(_08985_),
    .B2(_08996_),
    .X(_08997_));
 sky130_fd_sc_hd__a2bb2o_2 _23331_ (.A1_N(_08976_),
    .A2_N(_08997_),
    .B1(_08976_),
    .B2(_08997_),
    .X(_08998_));
 sky130_fd_sc_hd__a2bb2o_2 _23332_ (.A1_N(_08975_),
    .A2_N(_08998_),
    .B1(_08975_),
    .B2(_08998_),
    .X(_08999_));
 sky130_fd_sc_hd__o22a_2 _23333_ (.A1(_08901_),
    .A2(_08902_),
    .B1(_08896_),
    .B2(_08903_),
    .X(_09000_));
 sky130_fd_sc_hd__o22a_2 _23334_ (.A1(_08908_),
    .A2(_08914_),
    .B1(_08907_),
    .B2(_08915_),
    .X(_09001_));
 sky130_fd_sc_hd__o22a_2 _23335_ (.A1(_08559_),
    .A2(_06377_),
    .B1(_08431_),
    .B2(_06743_),
    .X(_09002_));
 sky130_fd_sc_hd__and4_2 _23336_ (.A(_08433_),
    .B(_06885_),
    .C(_11599_),
    .D(_11888_),
    .X(_09003_));
 sky130_fd_sc_hd__nor2_2 _23337_ (.A(_09002_),
    .B(_09003_),
    .Y(_09004_));
 sky130_fd_sc_hd__nor2_2 _23338_ (.A(_08437_),
    .B(_06625_),
    .Y(_09005_));
 sky130_fd_sc_hd__a2bb2o_2 _23339_ (.A1_N(_09004_),
    .A2_N(_09005_),
    .B1(_09004_),
    .B2(_09005_),
    .X(_09006_));
 sky130_fd_sc_hd__o22a_2 _23340_ (.A1(_08440_),
    .A2(_06904_),
    .B1(_08441_),
    .B2(_06754_),
    .X(_09007_));
 sky130_fd_sc_hd__and4_2 _23341_ (.A(_11586_),
    .B(_06499_),
    .C(_11590_),
    .D(_06627_),
    .X(_09008_));
 sky130_fd_sc_hd__nor2_2 _23342_ (.A(_09007_),
    .B(_09008_),
    .Y(_09009_));
 sky130_fd_sc_hd__nor2_2 _23343_ (.A(_05927_),
    .B(_06234_),
    .Y(_09010_));
 sky130_fd_sc_hd__a2bb2o_2 _23344_ (.A1_N(_09009_),
    .A2_N(_09010_),
    .B1(_09009_),
    .B2(_09010_),
    .X(_09011_));
 sky130_fd_sc_hd__a21oi_2 _23345_ (.A1(_08899_),
    .A2(_08900_),
    .B1(_08898_),
    .Y(_09012_));
 sky130_fd_sc_hd__a2bb2o_2 _23346_ (.A1_N(_09011_),
    .A2_N(_09012_),
    .B1(_09011_),
    .B2(_09012_),
    .X(_09013_));
 sky130_fd_sc_hd__a2bb2o_2 _23347_ (.A1_N(_09006_),
    .A2_N(_09013_),
    .B1(_09006_),
    .B2(_09013_),
    .X(_09014_));
 sky130_fd_sc_hd__a2bb2o_2 _23348_ (.A1_N(_09001_),
    .A2_N(_09014_),
    .B1(_09001_),
    .B2(_09014_),
    .X(_09015_));
 sky130_fd_sc_hd__a2bb2o_2 _23349_ (.A1_N(_09000_),
    .A2_N(_09015_),
    .B1(_09000_),
    .B2(_09015_),
    .X(_09016_));
 sky130_fd_sc_hd__a21oi_2 _23350_ (.A1(_08912_),
    .A2(_08913_),
    .B1(_08911_),
    .Y(_09017_));
 sky130_fd_sc_hd__a21oi_2 _23351_ (.A1(_08920_),
    .A2(_08921_),
    .B1(_08919_),
    .Y(_09018_));
 sky130_fd_sc_hd__o22a_2 _23352_ (.A1(_08909_),
    .A2(_07196_),
    .B1(_06442_),
    .B2(_05884_),
    .X(_09019_));
 sky130_fd_sc_hd__and4_2 _23353_ (.A(_11575_),
    .B(_06117_),
    .C(_08456_),
    .D(_11905_),
    .X(_09020_));
 sky130_fd_sc_hd__nor2_2 _23354_ (.A(_09019_),
    .B(_09020_),
    .Y(_09021_));
 sky130_fd_sc_hd__nor2_2 _23355_ (.A(_06273_),
    .B(_05893_),
    .Y(_09022_));
 sky130_fd_sc_hd__a2bb2o_2 _23356_ (.A1_N(_09021_),
    .A2_N(_09022_),
    .B1(_09021_),
    .B2(_09022_),
    .X(_09023_));
 sky130_fd_sc_hd__a2bb2o_2 _23357_ (.A1_N(_09018_),
    .A2_N(_09023_),
    .B1(_09018_),
    .B2(_09023_),
    .X(_09024_));
 sky130_fd_sc_hd__a2bb2o_2 _23358_ (.A1_N(_09017_),
    .A2_N(_09024_),
    .B1(_09017_),
    .B2(_09024_),
    .X(_09025_));
 sky130_fd_sc_hd__o22a_2 _23359_ (.A1(_08584_),
    .A2(_05429_),
    .B1(_06830_),
    .B2(_05895_),
    .X(_09026_));
 sky130_fd_sc_hd__and4_2 _23360_ (.A(_11567_),
    .B(_11915_),
    .C(_11571_),
    .D(_11913_),
    .X(_09027_));
 sky130_fd_sc_hd__nor2_2 _23361_ (.A(_09026_),
    .B(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__nor2_2 _23362_ (.A(_06687_),
    .B(_05704_),
    .Y(_09029_));
 sky130_fd_sc_hd__a2bb2o_2 _23363_ (.A1_N(_09028_),
    .A2_N(_09029_),
    .B1(_09028_),
    .B2(_09029_),
    .X(_09030_));
 sky130_fd_sc_hd__or2_2 _23364_ (.A(_08098_),
    .B(_05420_),
    .X(_09031_));
 sky130_fd_sc_hd__and4_2 _23365_ (.A(_07686_),
    .B(_05168_),
    .C(_08100_),
    .D(_11919_),
    .X(_09032_));
 sky130_fd_sc_hd__o22a_2 _23366_ (.A1(_08592_),
    .A2(_11922_),
    .B1(_07545_),
    .B2(_05255_),
    .X(_09033_));
 sky130_fd_sc_hd__or2_2 _23367_ (.A(_09032_),
    .B(_09033_),
    .X(_09034_));
 sky130_fd_sc_hd__a2bb2o_2 _23368_ (.A1_N(_09031_),
    .A2_N(_09034_),
    .B1(_09031_),
    .B2(_09034_),
    .X(_09035_));
 sky130_fd_sc_hd__o21ba_2 _23369_ (.A1(_08923_),
    .A2(_08926_),
    .B1_N(_08924_),
    .X(_09036_));
 sky130_fd_sc_hd__a2bb2o_2 _23370_ (.A1_N(_09035_),
    .A2_N(_09036_),
    .B1(_09035_),
    .B2(_09036_),
    .X(_09037_));
 sky130_fd_sc_hd__a2bb2o_2 _23371_ (.A1_N(_09030_),
    .A2_N(_09037_),
    .B1(_09030_),
    .B2(_09037_),
    .X(_09038_));
 sky130_fd_sc_hd__o22a_2 _23372_ (.A1(_08927_),
    .A2(_08928_),
    .B1(_08922_),
    .B2(_08929_),
    .X(_09039_));
 sky130_fd_sc_hd__a2bb2o_2 _23373_ (.A1_N(_09038_),
    .A2_N(_09039_),
    .B1(_09038_),
    .B2(_09039_),
    .X(_09040_));
 sky130_fd_sc_hd__a2bb2o_2 _23374_ (.A1_N(_09025_),
    .A2_N(_09040_),
    .B1(_09025_),
    .B2(_09040_),
    .X(_09041_));
 sky130_fd_sc_hd__o22a_2 _23375_ (.A1(_08930_),
    .A2(_08931_),
    .B1(_08916_),
    .B2(_08932_),
    .X(_09042_));
 sky130_fd_sc_hd__a2bb2o_2 _23376_ (.A1_N(_09041_),
    .A2_N(_09042_),
    .B1(_09041_),
    .B2(_09042_),
    .X(_09043_));
 sky130_fd_sc_hd__a2bb2o_2 _23377_ (.A1_N(_09016_),
    .A2_N(_09043_),
    .B1(_09016_),
    .B2(_09043_),
    .X(_09044_));
 sky130_fd_sc_hd__o22a_2 _23378_ (.A1(_08933_),
    .A2(_08934_),
    .B1(_08906_),
    .B2(_08935_),
    .X(_09045_));
 sky130_fd_sc_hd__a2bb2o_2 _23379_ (.A1_N(_09044_),
    .A2_N(_09045_),
    .B1(_09044_),
    .B2(_09045_),
    .X(_09046_));
 sky130_fd_sc_hd__a2bb2o_2 _23380_ (.A1_N(_08999_),
    .A2_N(_09046_),
    .B1(_08999_),
    .B2(_09046_),
    .X(_09047_));
 sky130_fd_sc_hd__o22a_2 _23381_ (.A1(_08936_),
    .A2(_08937_),
    .B1(_08889_),
    .B2(_08938_),
    .X(_09048_));
 sky130_fd_sc_hd__a2bb2o_2 _23382_ (.A1_N(_09047_),
    .A2_N(_09048_),
    .B1(_09047_),
    .B2(_09048_),
    .X(_09049_));
 sky130_fd_sc_hd__a2bb2o_2 _23383_ (.A1_N(_08974_),
    .A2_N(_09049_),
    .B1(_08974_),
    .B2(_09049_),
    .X(_09050_));
 sky130_fd_sc_hd__o22a_2 _23384_ (.A1(_08939_),
    .A2(_08940_),
    .B1(_08863_),
    .B2(_08941_),
    .X(_09051_));
 sky130_fd_sc_hd__a2bb2o_2 _23385_ (.A1_N(_09050_),
    .A2_N(_09051_),
    .B1(_09050_),
    .B2(_09051_),
    .X(_09052_));
 sky130_fd_sc_hd__a2bb2o_2 _23386_ (.A1_N(_08961_),
    .A2_N(_09052_),
    .B1(_08961_),
    .B2(_09052_),
    .X(_09053_));
 sky130_fd_sc_hd__o22a_2 _23387_ (.A1(_08942_),
    .A2(_08943_),
    .B1(_08845_),
    .B2(_08944_),
    .X(_09054_));
 sky130_fd_sc_hd__a2bb2o_2 _23388_ (.A1_N(_09053_),
    .A2_N(_09054_),
    .B1(_09053_),
    .B2(_09054_),
    .X(_09055_));
 sky130_fd_sc_hd__a2bb2o_2 _23389_ (.A1_N(_08844_),
    .A2_N(_09055_),
    .B1(_08844_),
    .B2(_09055_),
    .X(_09056_));
 sky130_fd_sc_hd__or2_2 _23390_ (.A(_08958_),
    .B(_09056_),
    .X(_09057_));
 sky130_fd_sc_hd__a21bo_2 _23391_ (.A1(_08958_),
    .A2(_09056_),
    .B1_N(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__o21ai_2 _23392_ (.A1(_08951_),
    .A2(_08956_),
    .B1(_08950_),
    .Y(_09059_));
 sky130_fd_sc_hd__a2bb2o_2 _23393_ (.A1_N(_09058_),
    .A2_N(_09059_),
    .B1(_09058_),
    .B2(_09059_),
    .X(_02664_));
 sky130_fd_sc_hd__o22a_2 _23394_ (.A1(_08963_),
    .A2(_08972_),
    .B1(_08962_),
    .B2(_08973_),
    .X(_09060_));
 sky130_fd_sc_hd__or2_2 _23395_ (.A(_08373_),
    .B(_09060_),
    .X(_09061_));
 sky130_fd_sc_hd__a21bo_2 _23396_ (.A1(_08375_),
    .A2(_09060_),
    .B1_N(_09061_),
    .X(_09062_));
 sky130_fd_sc_hd__o22a_2 _23397_ (.A1(_08968_),
    .A2(_08969_),
    .B1(_08623_),
    .B2(_08971_),
    .X(_09063_));
 sky130_fd_sc_hd__o22a_2 _23398_ (.A1(_08976_),
    .A2(_08997_),
    .B1(_08975_),
    .B2(_08998_),
    .X(_09064_));
 sky130_fd_sc_hd__o22a_2 _23399_ (.A1(_08978_),
    .A2(_08983_),
    .B1(_08757_),
    .B2(_08984_),
    .X(_09065_));
 sky130_fd_sc_hd__a2bb2o_2 _23400_ (.A1_N(_08853_),
    .A2_N(_09065_),
    .B1(_08853_),
    .B2(_09065_),
    .X(_09066_));
 sky130_fd_sc_hd__a2bb2o_2 _23401_ (.A1_N(_08966_),
    .A2_N(_09066_),
    .B1(_08966_),
    .B2(_09066_),
    .X(_09067_));
 sky130_fd_sc_hd__o22a_2 _23402_ (.A1(_08853_),
    .A2(_08964_),
    .B1(_08965_),
    .B2(_08966_),
    .X(_09068_));
 sky130_fd_sc_hd__o2bb2ai_2 _23403_ (.A1_N(_09067_),
    .A2_N(_09068_),
    .B1(_09067_),
    .B2(_09068_),
    .Y(_09069_));
 sky130_fd_sc_hd__a2bb2o_2 _23404_ (.A1_N(_08378_),
    .A2_N(_09069_),
    .B1(_08378_),
    .B2(_09069_),
    .X(_09070_));
 sky130_fd_sc_hd__a2bb2o_2 _23405_ (.A1_N(_09064_),
    .A2_N(_09070_),
    .B1(_09064_),
    .B2(_09070_),
    .X(_09071_));
 sky130_fd_sc_hd__a2bb2o_2 _23406_ (.A1_N(_09063_),
    .A2_N(_09071_),
    .B1(_09063_),
    .B2(_09071_),
    .X(_09072_));
 sky130_fd_sc_hd__o22a_2 _23407_ (.A1(_08994_),
    .A2(_08995_),
    .B1(_08985_),
    .B2(_08996_),
    .X(_09073_));
 sky130_fd_sc_hd__o22a_2 _23408_ (.A1(_09001_),
    .A2(_09014_),
    .B1(_09000_),
    .B2(_09015_),
    .X(_09074_));
 sky130_fd_sc_hd__buf_1 _23409_ (.A(_08757_),
    .X(_09075_));
 sky130_fd_sc_hd__or4_2 _23410_ (.A(_10587_),
    .B(_05132_),
    .C(_10587_),
    .D(_07626_),
    .X(_09076_));
 sky130_fd_sc_hd__a22o_2 _23411_ (.A1(_07870_),
    .A2(_11611_),
    .B1(_07870_),
    .B2(_11608_),
    .X(_09077_));
 sky130_fd_sc_hd__nand2_2 _23412_ (.A(_09076_),
    .B(_09077_),
    .Y(_09078_));
 sky130_fd_sc_hd__o22a_2 _23413_ (.A1(_08869_),
    .A2(_08980_),
    .B1(_05057_),
    .B2(_08979_),
    .X(_09079_));
 sky130_fd_sc_hd__a2bb2oi_2 _23414_ (.A1_N(_09078_),
    .A2_N(_09079_),
    .B1(_09078_),
    .B2(_09079_),
    .Y(_09080_));
 sky130_fd_sc_hd__a2bb2o_2 _23415_ (.A1_N(_09075_),
    .A2_N(_09080_),
    .B1(_09075_),
    .B2(_09080_),
    .X(_09081_));
 sky130_fd_sc_hd__a21oi_2 _23416_ (.A1(_08990_),
    .A2(_08991_),
    .B1(_08989_),
    .Y(_09082_));
 sky130_fd_sc_hd__a21oi_2 _23417_ (.A1(_09004_),
    .A2(_09005_),
    .B1(_09003_),
    .Y(_09083_));
 sky130_fd_sc_hd__o22a_2 _23418_ (.A1(_07918_),
    .A2(_07009_),
    .B1(_05389_),
    .B2(_07023_),
    .X(_09084_));
 sky130_fd_sc_hd__and4_2 _23419_ (.A(_11603_),
    .B(_07587_),
    .C(_11606_),
    .D(_11876_),
    .X(_09085_));
 sky130_fd_sc_hd__nor2_2 _23420_ (.A(_09084_),
    .B(_09085_),
    .Y(_09086_));
 sky130_fd_sc_hd__nor2_2 _23421_ (.A(_05310_),
    .B(_07160_),
    .Y(_09087_));
 sky130_fd_sc_hd__a2bb2o_2 _23422_ (.A1_N(_09086_),
    .A2_N(_09087_),
    .B1(_09086_),
    .B2(_09087_),
    .X(_09088_));
 sky130_fd_sc_hd__a2bb2o_2 _23423_ (.A1_N(_09083_),
    .A2_N(_09088_),
    .B1(_09083_),
    .B2(_09088_),
    .X(_09089_));
 sky130_fd_sc_hd__a2bb2o_2 _23424_ (.A1_N(_09082_),
    .A2_N(_09089_),
    .B1(_09082_),
    .B2(_09089_),
    .X(_09090_));
 sky130_fd_sc_hd__o22a_2 _23425_ (.A1(_08987_),
    .A2(_08992_),
    .B1(_08986_),
    .B2(_08993_),
    .X(_09091_));
 sky130_fd_sc_hd__a2bb2o_2 _23426_ (.A1_N(_09090_),
    .A2_N(_09091_),
    .B1(_09090_),
    .B2(_09091_),
    .X(_09092_));
 sky130_fd_sc_hd__a2bb2o_2 _23427_ (.A1_N(_09081_),
    .A2_N(_09092_),
    .B1(_09081_),
    .B2(_09092_),
    .X(_09093_));
 sky130_fd_sc_hd__a2bb2o_2 _23428_ (.A1_N(_09074_),
    .A2_N(_09093_),
    .B1(_09074_),
    .B2(_09093_),
    .X(_09094_));
 sky130_fd_sc_hd__a2bb2o_2 _23429_ (.A1_N(_09073_),
    .A2_N(_09094_),
    .B1(_09073_),
    .B2(_09094_),
    .X(_09095_));
 sky130_fd_sc_hd__o22a_2 _23430_ (.A1(_09011_),
    .A2(_09012_),
    .B1(_09006_),
    .B2(_09013_),
    .X(_09096_));
 sky130_fd_sc_hd__o22a_2 _23431_ (.A1(_09018_),
    .A2(_09023_),
    .B1(_09017_),
    .B2(_09024_),
    .X(_09097_));
 sky130_fd_sc_hd__o22a_2 _23432_ (.A1(_08559_),
    .A2(_06496_),
    .B1(_05660_),
    .B2(_06879_),
    .X(_09098_));
 sky130_fd_sc_hd__and4_2 _23433_ (.A(_11594_),
    .B(_11888_),
    .C(_11599_),
    .D(_07155_),
    .X(_09099_));
 sky130_fd_sc_hd__nor2_2 _23434_ (.A(_09098_),
    .B(_09099_),
    .Y(_09100_));
 sky130_fd_sc_hd__nor2_2 _23435_ (.A(_05563_),
    .B(_07008_),
    .Y(_09101_));
 sky130_fd_sc_hd__a2bb2o_2 _23436_ (.A1_N(_09100_),
    .A2_N(_09101_),
    .B1(_09100_),
    .B2(_09101_),
    .X(_09102_));
 sky130_fd_sc_hd__buf_1 _23437_ (.A(_06818_),
    .X(_09103_));
 sky130_fd_sc_hd__o22a_2 _23438_ (.A1(_09103_),
    .A2(_06754_),
    .B1(_08441_),
    .B2(_06233_),
    .X(_09104_));
 sky130_fd_sc_hd__and4_2 _23439_ (.A(_11586_),
    .B(_06627_),
    .C(_11590_),
    .D(_06752_),
    .X(_09105_));
 sky130_fd_sc_hd__nor2_2 _23440_ (.A(_09104_),
    .B(_09105_),
    .Y(_09106_));
 sky130_fd_sc_hd__nor2_2 _23441_ (.A(_05927_),
    .B(_06617_),
    .Y(_09107_));
 sky130_fd_sc_hd__a2bb2o_2 _23442_ (.A1_N(_09106_),
    .A2_N(_09107_),
    .B1(_09106_),
    .B2(_09107_),
    .X(_09108_));
 sky130_fd_sc_hd__a21oi_2 _23443_ (.A1(_09009_),
    .A2(_09010_),
    .B1(_09008_),
    .Y(_09109_));
 sky130_fd_sc_hd__a2bb2o_2 _23444_ (.A1_N(_09108_),
    .A2_N(_09109_),
    .B1(_09108_),
    .B2(_09109_),
    .X(_09110_));
 sky130_fd_sc_hd__a2bb2o_2 _23445_ (.A1_N(_09102_),
    .A2_N(_09110_),
    .B1(_09102_),
    .B2(_09110_),
    .X(_09111_));
 sky130_fd_sc_hd__a2bb2o_2 _23446_ (.A1_N(_09097_),
    .A2_N(_09111_),
    .B1(_09097_),
    .B2(_09111_),
    .X(_09112_));
 sky130_fd_sc_hd__a2bb2o_2 _23447_ (.A1_N(_09096_),
    .A2_N(_09112_),
    .B1(_09096_),
    .B2(_09112_),
    .X(_09113_));
 sky130_fd_sc_hd__a21oi_2 _23448_ (.A1(_09021_),
    .A2(_09022_),
    .B1(_09020_),
    .Y(_09114_));
 sky130_fd_sc_hd__a21oi_2 _23449_ (.A1(_09028_),
    .A2(_09029_),
    .B1(_09027_),
    .Y(_09115_));
 sky130_fd_sc_hd__o22a_2 _23450_ (.A1(_08909_),
    .A2(_05884_),
    .B1(_06442_),
    .B2(_05892_),
    .X(_09116_));
 sky130_fd_sc_hd__and4_2 _23451_ (.A(_11575_),
    .B(_06240_),
    .C(_08456_),
    .D(_11902_),
    .X(_09117_));
 sky130_fd_sc_hd__nor2_2 _23452_ (.A(_09116_),
    .B(_09117_),
    .Y(_09118_));
 sky130_fd_sc_hd__nor2_2 _23453_ (.A(_06273_),
    .B(_08057_),
    .Y(_09119_));
 sky130_fd_sc_hd__a2bb2o_2 _23454_ (.A1_N(_09118_),
    .A2_N(_09119_),
    .B1(_09118_),
    .B2(_09119_),
    .X(_09120_));
 sky130_fd_sc_hd__a2bb2o_2 _23455_ (.A1_N(_09115_),
    .A2_N(_09120_),
    .B1(_09115_),
    .B2(_09120_),
    .X(_09121_));
 sky130_fd_sc_hd__a2bb2o_2 _23456_ (.A1_N(_09114_),
    .A2_N(_09121_),
    .B1(_09114_),
    .B2(_09121_),
    .X(_09122_));
 sky130_fd_sc_hd__o22a_2 _23457_ (.A1(_08584_),
    .A2(_05895_),
    .B1(_06833_),
    .B2(_05607_),
    .X(_09123_));
 sky130_fd_sc_hd__and4_2 _23458_ (.A(_07680_),
    .B(_05897_),
    .C(_11571_),
    .D(_11911_),
    .X(_09124_));
 sky130_fd_sc_hd__nor2_2 _23459_ (.A(_09123_),
    .B(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__nor2_2 _23460_ (.A(_07822_),
    .B(_05816_),
    .Y(_09126_));
 sky130_fd_sc_hd__a2bb2o_2 _23461_ (.A1_N(_09125_),
    .A2_N(_09126_),
    .B1(_09125_),
    .B2(_09126_),
    .X(_09127_));
 sky130_fd_sc_hd__buf_1 _23462_ (.A(_07393_),
    .X(_09128_));
 sky130_fd_sc_hd__and4_2 _23463_ (.A(_09128_),
    .B(_05255_),
    .C(_11560_),
    .D(_11916_),
    .X(_09129_));
 sky130_fd_sc_hd__o22a_2 _23464_ (.A1(_10597_),
    .A2(_11919_),
    .B1(_07247_),
    .B2(_05342_),
    .X(_09130_));
 sky130_fd_sc_hd__nor2_2 _23465_ (.A(_09129_),
    .B(_09130_),
    .Y(_09131_));
 sky130_fd_sc_hd__nor2_2 _23466_ (.A(_07828_),
    .B(_06134_),
    .Y(_09132_));
 sky130_fd_sc_hd__a2bb2o_2 _23467_ (.A1_N(_09131_),
    .A2_N(_09132_),
    .B1(_09131_),
    .B2(_09132_),
    .X(_09133_));
 sky130_fd_sc_hd__o21ba_2 _23468_ (.A1(_09031_),
    .A2(_09034_),
    .B1_N(_09032_),
    .X(_09134_));
 sky130_fd_sc_hd__a2bb2o_2 _23469_ (.A1_N(_09133_),
    .A2_N(_09134_),
    .B1(_09133_),
    .B2(_09134_),
    .X(_09135_));
 sky130_fd_sc_hd__a2bb2o_2 _23470_ (.A1_N(_09127_),
    .A2_N(_09135_),
    .B1(_09127_),
    .B2(_09135_),
    .X(_09136_));
 sky130_fd_sc_hd__o22a_2 _23471_ (.A1(_09035_),
    .A2(_09036_),
    .B1(_09030_),
    .B2(_09037_),
    .X(_09137_));
 sky130_fd_sc_hd__a2bb2o_2 _23472_ (.A1_N(_09136_),
    .A2_N(_09137_),
    .B1(_09136_),
    .B2(_09137_),
    .X(_09138_));
 sky130_fd_sc_hd__a2bb2o_2 _23473_ (.A1_N(_09122_),
    .A2_N(_09138_),
    .B1(_09122_),
    .B2(_09138_),
    .X(_09139_));
 sky130_fd_sc_hd__o22a_2 _23474_ (.A1(_09038_),
    .A2(_09039_),
    .B1(_09025_),
    .B2(_09040_),
    .X(_09140_));
 sky130_fd_sc_hd__a2bb2o_2 _23475_ (.A1_N(_09139_),
    .A2_N(_09140_),
    .B1(_09139_),
    .B2(_09140_),
    .X(_09141_));
 sky130_fd_sc_hd__a2bb2o_2 _23476_ (.A1_N(_09113_),
    .A2_N(_09141_),
    .B1(_09113_),
    .B2(_09141_),
    .X(_09142_));
 sky130_fd_sc_hd__o22a_2 _23477_ (.A1(_09041_),
    .A2(_09042_),
    .B1(_09016_),
    .B2(_09043_),
    .X(_09143_));
 sky130_fd_sc_hd__a2bb2o_2 _23478_ (.A1_N(_09142_),
    .A2_N(_09143_),
    .B1(_09142_),
    .B2(_09143_),
    .X(_09144_));
 sky130_fd_sc_hd__a2bb2o_2 _23479_ (.A1_N(_09095_),
    .A2_N(_09144_),
    .B1(_09095_),
    .B2(_09144_),
    .X(_09145_));
 sky130_fd_sc_hd__o22a_2 _23480_ (.A1(_09044_),
    .A2(_09045_),
    .B1(_08999_),
    .B2(_09046_),
    .X(_09146_));
 sky130_fd_sc_hd__a2bb2o_2 _23481_ (.A1_N(_09145_),
    .A2_N(_09146_),
    .B1(_09145_),
    .B2(_09146_),
    .X(_09147_));
 sky130_fd_sc_hd__a2bb2o_2 _23482_ (.A1_N(_09072_),
    .A2_N(_09147_),
    .B1(_09072_),
    .B2(_09147_),
    .X(_09148_));
 sky130_fd_sc_hd__o22a_2 _23483_ (.A1(_09047_),
    .A2(_09048_),
    .B1(_08974_),
    .B2(_09049_),
    .X(_09149_));
 sky130_fd_sc_hd__a2bb2o_2 _23484_ (.A1_N(_09148_),
    .A2_N(_09149_),
    .B1(_09148_),
    .B2(_09149_),
    .X(_09150_));
 sky130_fd_sc_hd__a2bb2o_2 _23485_ (.A1_N(_09062_),
    .A2_N(_09150_),
    .B1(_09062_),
    .B2(_09150_),
    .X(_09151_));
 sky130_fd_sc_hd__o22a_2 _23486_ (.A1(_09050_),
    .A2(_09051_),
    .B1(_08961_),
    .B2(_09052_),
    .X(_09152_));
 sky130_fd_sc_hd__a2bb2o_2 _23487_ (.A1_N(_09151_),
    .A2_N(_09152_),
    .B1(_09151_),
    .B2(_09152_),
    .X(_09153_));
 sky130_fd_sc_hd__a2bb2o_2 _23488_ (.A1_N(_08960_),
    .A2_N(_09153_),
    .B1(_08960_),
    .B2(_09153_),
    .X(_09154_));
 sky130_fd_sc_hd__o22a_2 _23489_ (.A1(_09053_),
    .A2(_09054_),
    .B1(_08844_),
    .B2(_09055_),
    .X(_09155_));
 sky130_fd_sc_hd__or2_2 _23490_ (.A(_09154_),
    .B(_09155_),
    .X(_09156_));
 sky130_fd_sc_hd__a21bo_2 _23491_ (.A1(_09154_),
    .A2(_09155_),
    .B1_N(_09156_),
    .X(_09157_));
 sky130_fd_sc_hd__a22o_2 _23492_ (.A1(_08958_),
    .A2(_09056_),
    .B1(_08950_),
    .B2(_09057_),
    .X(_09158_));
 sky130_fd_sc_hd__o31a_2 _23493_ (.A1(_08951_),
    .A2(_09058_),
    .A3(_08956_),
    .B1(_09158_),
    .X(_09159_));
 sky130_fd_sc_hd__a2bb2oi_2 _23494_ (.A1_N(_09157_),
    .A2_N(_09159_),
    .B1(_09157_),
    .B2(_09159_),
    .Y(_02665_));
 sky130_fd_sc_hd__o22a_2 _23495_ (.A1(_09151_),
    .A2(_09152_),
    .B1(_08960_),
    .B2(_09153_),
    .X(_09160_));
 sky130_fd_sc_hd__o22a_2 _23496_ (.A1(_09064_),
    .A2(_09070_),
    .B1(_09063_),
    .B2(_09071_),
    .X(_09161_));
 sky130_fd_sc_hd__or2_2 _23497_ (.A(_08373_),
    .B(_09161_),
    .X(_09162_));
 sky130_fd_sc_hd__a21bo_2 _23498_ (.A1(_08374_),
    .A2(_09161_),
    .B1_N(_09162_),
    .X(_09163_));
 sky130_fd_sc_hd__o22a_2 _23499_ (.A1(_09067_),
    .A2(_09068_),
    .B1(_08379_),
    .B2(_09069_),
    .X(_09164_));
 sky130_fd_sc_hd__o22a_2 _23500_ (.A1(_09074_),
    .A2(_09093_),
    .B1(_09073_),
    .B2(_09094_),
    .X(_09165_));
 sky130_fd_sc_hd__o22a_2 _23501_ (.A1(_08853_),
    .A2(_09065_),
    .B1(_08966_),
    .B2(_09066_),
    .X(_09166_));
 sky130_fd_sc_hd__o22ai_2 _23502_ (.A1(_09075_),
    .A2(_09080_),
    .B1(_05057_),
    .B2(_09076_),
    .Y(_09167_));
 sky130_fd_sc_hd__and3_2 _23503_ (.A(_08389_),
    .B(_08849_),
    .C(_08627_),
    .X(_09168_));
 sky130_fd_sc_hd__o21ba_2 _23504_ (.A1(_08743_),
    .A2(_08850_),
    .B1_N(_09168_),
    .X(_09169_));
 sky130_fd_sc_hd__a2bb2o_2 _23505_ (.A1_N(_09167_),
    .A2_N(_09169_),
    .B1(_09167_),
    .B2(_09169_),
    .X(_09170_));
 sky130_fd_sc_hd__o2bb2ai_2 _23506_ (.A1_N(_09166_),
    .A2_N(_09170_),
    .B1(_09166_),
    .B2(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__a2bb2o_2 _23507_ (.A1_N(_08623_),
    .A2_N(_09171_),
    .B1(_08623_),
    .B2(_09171_),
    .X(_09172_));
 sky130_fd_sc_hd__a2bb2o_2 _23508_ (.A1_N(_09165_),
    .A2_N(_09172_),
    .B1(_09165_),
    .B2(_09172_),
    .X(_09173_));
 sky130_fd_sc_hd__a2bb2o_2 _23509_ (.A1_N(_09164_),
    .A2_N(_09173_),
    .B1(_09164_),
    .B2(_09173_),
    .X(_09174_));
 sky130_fd_sc_hd__o22a_2 _23510_ (.A1(_09090_),
    .A2(_09091_),
    .B1(_09081_),
    .B2(_09092_),
    .X(_09175_));
 sky130_fd_sc_hd__o22a_2 _23511_ (.A1(_09097_),
    .A2(_09111_),
    .B1(_09096_),
    .B2(_09112_),
    .X(_09176_));
 sky130_fd_sc_hd__o22ai_2 _23512_ (.A1(_05057_),
    .A2(_09076_),
    .B1(_08869_),
    .B2(_09077_),
    .Y(_09177_));
 sky130_fd_sc_hd__a2bb2o_2 _23513_ (.A1_N(_09075_),
    .A2_N(_09177_),
    .B1(_09075_),
    .B2(_09177_),
    .X(_09178_));
 sky130_fd_sc_hd__a21oi_2 _23514_ (.A1(_09086_),
    .A2(_09087_),
    .B1(_09085_),
    .Y(_09179_));
 sky130_fd_sc_hd__a21oi_2 _23515_ (.A1(_09100_),
    .A2(_09101_),
    .B1(_09099_),
    .Y(_09180_));
 sky130_fd_sc_hd__o22a_2 _23516_ (.A1(_07918_),
    .A2(_07023_),
    .B1(_05389_),
    .B2(_07159_),
    .X(_09181_));
 sky130_fd_sc_hd__and4_2 _23517_ (.A(_11603_),
    .B(_11877_),
    .C(_11606_),
    .D(_11873_),
    .X(_09182_));
 sky130_fd_sc_hd__nor2_2 _23518_ (.A(_09181_),
    .B(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__or2_2 _23519_ (.A(_10586_),
    .B(_05393_),
    .X(_09184_));
 sky130_vsdinv _23520_ (.A(_09184_),
    .Y(_09185_));
 sky130_fd_sc_hd__a2bb2o_2 _23521_ (.A1_N(_09183_),
    .A2_N(_09185_),
    .B1(_09183_),
    .B2(_09185_),
    .X(_09186_));
 sky130_fd_sc_hd__a2bb2o_2 _23522_ (.A1_N(_09180_),
    .A2_N(_09186_),
    .B1(_09180_),
    .B2(_09186_),
    .X(_09187_));
 sky130_fd_sc_hd__a2bb2o_2 _23523_ (.A1_N(_09179_),
    .A2_N(_09187_),
    .B1(_09179_),
    .B2(_09187_),
    .X(_09188_));
 sky130_fd_sc_hd__o22a_2 _23524_ (.A1(_09083_),
    .A2(_09088_),
    .B1(_09082_),
    .B2(_09089_),
    .X(_09189_));
 sky130_fd_sc_hd__a2bb2o_2 _23525_ (.A1_N(_09188_),
    .A2_N(_09189_),
    .B1(_09188_),
    .B2(_09189_),
    .X(_09190_));
 sky130_fd_sc_hd__a2bb2o_2 _23526_ (.A1_N(_09178_),
    .A2_N(_09190_),
    .B1(_09178_),
    .B2(_09190_),
    .X(_09191_));
 sky130_fd_sc_hd__a2bb2o_2 _23527_ (.A1_N(_09176_),
    .A2_N(_09191_),
    .B1(_09176_),
    .B2(_09191_),
    .X(_09192_));
 sky130_fd_sc_hd__a2bb2o_2 _23528_ (.A1_N(_09175_),
    .A2_N(_09192_),
    .B1(_09175_),
    .B2(_09192_),
    .X(_09193_));
 sky130_fd_sc_hd__o22a_2 _23529_ (.A1(_09108_),
    .A2(_09109_),
    .B1(_09102_),
    .B2(_09110_),
    .X(_09194_));
 sky130_fd_sc_hd__o22a_2 _23530_ (.A1(_09115_),
    .A2(_09120_),
    .B1(_09114_),
    .B2(_09121_),
    .X(_09195_));
 sky130_fd_sc_hd__o22a_2 _23531_ (.A1(_08559_),
    .A2(_06624_),
    .B1(_08431_),
    .B2(_07007_),
    .X(_09196_));
 sky130_fd_sc_hd__and4_2 _23532_ (.A(_08433_),
    .B(_07155_),
    .C(_08434_),
    .D(_11882_),
    .X(_09197_));
 sky130_fd_sc_hd__nor2_2 _23533_ (.A(_09196_),
    .B(_09197_),
    .Y(_09198_));
 sky130_fd_sc_hd__nor2_2 _23534_ (.A(_05563_),
    .B(_07289_),
    .Y(_09199_));
 sky130_fd_sc_hd__a2bb2o_2 _23535_ (.A1_N(_09198_),
    .A2_N(_09199_),
    .B1(_09198_),
    .B2(_09199_),
    .X(_09200_));
 sky130_fd_sc_hd__o22a_2 _23536_ (.A1(_09103_),
    .A2(_06233_),
    .B1(_06031_),
    .B2(_06616_),
    .X(_09201_));
 sky130_fd_sc_hd__and4_2 _23537_ (.A(_11586_),
    .B(_06752_),
    .C(_11590_),
    .D(_06885_),
    .X(_09202_));
 sky130_fd_sc_hd__nor2_2 _23538_ (.A(_09201_),
    .B(_09202_),
    .Y(_09203_));
 sky130_fd_sc_hd__nor2_2 _23539_ (.A(_05927_),
    .B(_06497_),
    .Y(_09204_));
 sky130_fd_sc_hd__a2bb2o_2 _23540_ (.A1_N(_09203_),
    .A2_N(_09204_),
    .B1(_09203_),
    .B2(_09204_),
    .X(_09205_));
 sky130_fd_sc_hd__a21oi_2 _23541_ (.A1(_09106_),
    .A2(_09107_),
    .B1(_09105_),
    .Y(_09206_));
 sky130_fd_sc_hd__a2bb2o_2 _23542_ (.A1_N(_09205_),
    .A2_N(_09206_),
    .B1(_09205_),
    .B2(_09206_),
    .X(_09207_));
 sky130_fd_sc_hd__a2bb2o_2 _23543_ (.A1_N(_09200_),
    .A2_N(_09207_),
    .B1(_09200_),
    .B2(_09207_),
    .X(_09208_));
 sky130_fd_sc_hd__a2bb2o_2 _23544_ (.A1_N(_09195_),
    .A2_N(_09208_),
    .B1(_09195_),
    .B2(_09208_),
    .X(_09209_));
 sky130_fd_sc_hd__a2bb2o_2 _23545_ (.A1_N(_09194_),
    .A2_N(_09209_),
    .B1(_09194_),
    .B2(_09209_),
    .X(_09210_));
 sky130_fd_sc_hd__a21oi_2 _23546_ (.A1(_09118_),
    .A2(_09119_),
    .B1(_09117_),
    .Y(_09211_));
 sky130_fd_sc_hd__a21oi_2 _23547_ (.A1(_09125_),
    .A2(_09126_),
    .B1(_09124_),
    .Y(_09212_));
 sky130_fd_sc_hd__o22a_2 _23548_ (.A1(_08909_),
    .A2(_06501_),
    .B1(_06442_),
    .B2(_06502_),
    .X(_09213_));
 sky130_fd_sc_hd__and4_2 _23549_ (.A(_11575_),
    .B(_06372_),
    .C(_11581_),
    .D(_06499_),
    .X(_09214_));
 sky130_fd_sc_hd__nor2_2 _23550_ (.A(_09213_),
    .B(_09214_),
    .Y(_09215_));
 sky130_fd_sc_hd__nor2_2 _23551_ (.A(_06273_),
    .B(_06112_),
    .Y(_09216_));
 sky130_fd_sc_hd__a2bb2o_2 _23552_ (.A1_N(_09215_),
    .A2_N(_09216_),
    .B1(_09215_),
    .B2(_09216_),
    .X(_09217_));
 sky130_fd_sc_hd__a2bb2o_2 _23553_ (.A1_N(_09212_),
    .A2_N(_09217_),
    .B1(_09212_),
    .B2(_09217_),
    .X(_09218_));
 sky130_fd_sc_hd__a2bb2o_2 _23554_ (.A1_N(_09211_),
    .A2_N(_09218_),
    .B1(_09211_),
    .B2(_09218_),
    .X(_09219_));
 sky130_fd_sc_hd__and4_2 _23555_ (.A(_07393_),
    .B(_05341_),
    .C(_11559_),
    .D(\pcpi_mul.rs1[16] ),
    .X(_09220_));
 sky130_fd_sc_hd__o22a_2 _23556_ (.A1(_08592_),
    .A2(_11916_),
    .B1(_07545_),
    .B2(_05427_),
    .X(_09221_));
 sky130_fd_sc_hd__nor2_2 _23557_ (.A(_09220_),
    .B(_09221_),
    .Y(_09222_));
 sky130_fd_sc_hd__nor2_2 _23558_ (.A(_07100_),
    .B(_05598_),
    .Y(_09223_));
 sky130_fd_sc_hd__a2bb2o_2 _23559_ (.A1_N(_09222_),
    .A2_N(_09223_),
    .B1(_09222_),
    .B2(_09223_),
    .X(_09224_));
 sky130_fd_sc_hd__a21oi_2 _23560_ (.A1(_09131_),
    .A2(_09132_),
    .B1(_09129_),
    .Y(_09225_));
 sky130_fd_sc_hd__o2bb2a_2 _23561_ (.A1_N(_09224_),
    .A2_N(_09225_),
    .B1(_09224_),
    .B2(_09225_),
    .X(_09226_));
 sky130_vsdinv _23562_ (.A(_09226_),
    .Y(_09227_));
 sky130_fd_sc_hd__o22a_2 _23563_ (.A1(_08584_),
    .A2(_07059_),
    .B1(_06833_),
    .B2(_05715_),
    .X(_09228_));
 sky130_fd_sc_hd__and4_2 _23564_ (.A(_07680_),
    .B(_06393_),
    .C(_07681_),
    .D(_11908_),
    .X(_09229_));
 sky130_fd_sc_hd__nor2_2 _23565_ (.A(_09228_),
    .B(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__nor2_2 _23566_ (.A(_07822_),
    .B(_05824_),
    .Y(_09231_));
 sky130_fd_sc_hd__a2bb2o_2 _23567_ (.A1_N(_09230_),
    .A2_N(_09231_),
    .B1(_09230_),
    .B2(_09231_),
    .X(_09232_));
 sky130_vsdinv _23568_ (.A(_09232_),
    .Y(_09233_));
 sky130_fd_sc_hd__a22o_2 _23569_ (.A1(_09227_),
    .A2(_09232_),
    .B1(_09226_),
    .B2(_09233_),
    .X(_09234_));
 sky130_fd_sc_hd__o22a_2 _23570_ (.A1(_09133_),
    .A2(_09134_),
    .B1(_09127_),
    .B2(_09135_),
    .X(_09235_));
 sky130_fd_sc_hd__a2bb2o_2 _23571_ (.A1_N(_09234_),
    .A2_N(_09235_),
    .B1(_09234_),
    .B2(_09235_),
    .X(_09236_));
 sky130_fd_sc_hd__a2bb2o_2 _23572_ (.A1_N(_09219_),
    .A2_N(_09236_),
    .B1(_09219_),
    .B2(_09236_),
    .X(_09237_));
 sky130_fd_sc_hd__o22a_2 _23573_ (.A1(_09136_),
    .A2(_09137_),
    .B1(_09122_),
    .B2(_09138_),
    .X(_09238_));
 sky130_fd_sc_hd__a2bb2o_2 _23574_ (.A1_N(_09237_),
    .A2_N(_09238_),
    .B1(_09237_),
    .B2(_09238_),
    .X(_09239_));
 sky130_fd_sc_hd__a2bb2o_2 _23575_ (.A1_N(_09210_),
    .A2_N(_09239_),
    .B1(_09210_),
    .B2(_09239_),
    .X(_09240_));
 sky130_fd_sc_hd__o22a_2 _23576_ (.A1(_09139_),
    .A2(_09140_),
    .B1(_09113_),
    .B2(_09141_),
    .X(_09241_));
 sky130_fd_sc_hd__a2bb2o_2 _23577_ (.A1_N(_09240_),
    .A2_N(_09241_),
    .B1(_09240_),
    .B2(_09241_),
    .X(_09242_));
 sky130_fd_sc_hd__a2bb2o_2 _23578_ (.A1_N(_09193_),
    .A2_N(_09242_),
    .B1(_09193_),
    .B2(_09242_),
    .X(_09243_));
 sky130_fd_sc_hd__o22a_2 _23579_ (.A1(_09142_),
    .A2(_09143_),
    .B1(_09095_),
    .B2(_09144_),
    .X(_09244_));
 sky130_fd_sc_hd__a2bb2o_2 _23580_ (.A1_N(_09243_),
    .A2_N(_09244_),
    .B1(_09243_),
    .B2(_09244_),
    .X(_09245_));
 sky130_fd_sc_hd__a2bb2o_2 _23581_ (.A1_N(_09174_),
    .A2_N(_09245_),
    .B1(_09174_),
    .B2(_09245_),
    .X(_09246_));
 sky130_fd_sc_hd__o22a_2 _23582_ (.A1(_09145_),
    .A2(_09146_),
    .B1(_09072_),
    .B2(_09147_),
    .X(_09247_));
 sky130_fd_sc_hd__a2bb2o_2 _23583_ (.A1_N(_09246_),
    .A2_N(_09247_),
    .B1(_09246_),
    .B2(_09247_),
    .X(_09248_));
 sky130_fd_sc_hd__a2bb2o_2 _23584_ (.A1_N(_09163_),
    .A2_N(_09248_),
    .B1(_09163_),
    .B2(_09248_),
    .X(_09249_));
 sky130_fd_sc_hd__o22a_2 _23585_ (.A1(_09148_),
    .A2(_09149_),
    .B1(_09062_),
    .B2(_09150_),
    .X(_09250_));
 sky130_fd_sc_hd__a2bb2o_2 _23586_ (.A1_N(_09249_),
    .A2_N(_09250_),
    .B1(_09249_),
    .B2(_09250_),
    .X(_09251_));
 sky130_fd_sc_hd__a2bb2o_2 _23587_ (.A1_N(_09061_),
    .A2_N(_09251_),
    .B1(_09061_),
    .B2(_09251_),
    .X(_09252_));
 sky130_fd_sc_hd__and2_2 _23588_ (.A(_09160_),
    .B(_09252_),
    .X(_09253_));
 sky130_fd_sc_hd__or2_2 _23589_ (.A(_09160_),
    .B(_09252_),
    .X(_09254_));
 sky130_fd_sc_hd__or2b_2 _23590_ (.A(_09253_),
    .B_N(_09254_),
    .X(_09255_));
 sky130_fd_sc_hd__o21ai_2 _23591_ (.A1(_09157_),
    .A2(_09159_),
    .B1(_09156_),
    .Y(_09256_));
 sky130_fd_sc_hd__a2bb2o_2 _23592_ (.A1_N(_09255_),
    .A2_N(_09256_),
    .B1(_09255_),
    .B2(_09256_),
    .X(_02666_));
 sky130_fd_sc_hd__buf_1 _23593_ (.A(_08842_),
    .X(_09257_));
 sky130_fd_sc_hd__buf_1 _23594_ (.A(_09257_),
    .X(_09258_));
 sky130_fd_sc_hd__o22a_2 _23595_ (.A1(_09165_),
    .A2(_09172_),
    .B1(_09164_),
    .B2(_09173_),
    .X(_09259_));
 sky130_fd_sc_hd__or2_2 _23596_ (.A(_09257_),
    .B(_09259_),
    .X(_09260_));
 sky130_fd_sc_hd__a21bo_2 _23597_ (.A1(_09258_),
    .A2(_09259_),
    .B1_N(_09260_),
    .X(_09261_));
 sky130_fd_sc_hd__buf_1 _23598_ (.A(_08379_),
    .X(_09262_));
 sky130_fd_sc_hd__o22a_2 _23599_ (.A1(_09166_),
    .A2(_09170_),
    .B1(_09262_),
    .B2(_09171_),
    .X(_09263_));
 sky130_fd_sc_hd__o22a_2 _23600_ (.A1(_09176_),
    .A2(_09191_),
    .B1(_09175_),
    .B2(_09192_),
    .X(_09264_));
 sky130_fd_sc_hd__o22a_2 _23601_ (.A1(_05057_),
    .A2(_09076_),
    .B1(_09075_),
    .B2(_09177_),
    .X(_09265_));
 sky130_fd_sc_hd__o22ai_2 _23602_ (.A1(_08743_),
    .A2(_08850_),
    .B1(_09167_),
    .B2(_09168_),
    .Y(_09266_));
 sky130_fd_sc_hd__o2bb2a_2 _23603_ (.A1_N(_09265_),
    .A2_N(_09266_),
    .B1(_09265_),
    .B2(_09266_),
    .X(_09267_));
 sky130_fd_sc_hd__a2bb2o_2 _23604_ (.A1_N(_09262_),
    .A2_N(_09267_),
    .B1(_09262_),
    .B2(_09267_),
    .X(_09268_));
 sky130_fd_sc_hd__a2bb2o_2 _23605_ (.A1_N(_09264_),
    .A2_N(_09268_),
    .B1(_09264_),
    .B2(_09268_),
    .X(_09269_));
 sky130_fd_sc_hd__a2bb2o_2 _23606_ (.A1_N(_09263_),
    .A2_N(_09269_),
    .B1(_09263_),
    .B2(_09269_),
    .X(_09270_));
 sky130_fd_sc_hd__buf_1 _23607_ (.A(_09178_),
    .X(_09271_));
 sky130_fd_sc_hd__buf_1 _23608_ (.A(_09271_),
    .X(_09272_));
 sky130_fd_sc_hd__o22a_2 _23609_ (.A1(_09188_),
    .A2(_09189_),
    .B1(_09272_),
    .B2(_09190_),
    .X(_09273_));
 sky130_fd_sc_hd__o22a_2 _23610_ (.A1(_09195_),
    .A2(_09208_),
    .B1(_09194_),
    .B2(_09209_),
    .X(_09274_));
 sky130_fd_sc_hd__a31o_2 _23611_ (.A1(\pcpi_mul.rs2[18] ),
    .A2(_07012_),
    .A3(_09198_),
    .B1(_09197_),
    .X(_09275_));
 sky130_fd_sc_hd__o22a_2 _23612_ (.A1(_07340_),
    .A2(_07732_),
    .B1(_07727_),
    .B2(_05392_),
    .X(_09276_));
 sky130_fd_sc_hd__and4_2 _23613_ (.A(_07342_),
    .B(_11873_),
    .C(_07868_),
    .D(_07343_),
    .X(_09277_));
 sky130_fd_sc_hd__or2_2 _23614_ (.A(_09276_),
    .B(_09277_),
    .X(_09278_));
 sky130_vsdinv _23615_ (.A(_09278_),
    .Y(_09279_));
 sky130_fd_sc_hd__o22a_2 _23616_ (.A1(_09184_),
    .A2(_09278_),
    .B1(_09185_),
    .B2(_09279_),
    .X(_09280_));
 sky130_vsdinv _23617_ (.A(_09275_),
    .Y(_09281_));
 sky130_vsdinv _23618_ (.A(_09280_),
    .Y(_09282_));
 sky130_fd_sc_hd__o22a_2 _23619_ (.A1(_09275_),
    .A2(_09280_),
    .B1(_09281_),
    .B2(_09282_),
    .X(_09283_));
 sky130_fd_sc_hd__buf_1 _23620_ (.A(_07870_),
    .X(_09284_));
 sky130_fd_sc_hd__a31o_2 _23621_ (.A1(_09284_),
    .A2(\pcpi_mul.rs2[15] ),
    .A3(_09183_),
    .B1(_09182_),
    .X(_09285_));
 sky130_vsdinv _23622_ (.A(_09283_),
    .Y(_09286_));
 sky130_vsdinv _23623_ (.A(_09285_),
    .Y(_09287_));
 sky130_fd_sc_hd__o22a_2 _23624_ (.A1(_09283_),
    .A2(_09285_),
    .B1(_09286_),
    .B2(_09287_),
    .X(_09288_));
 sky130_vsdinv _23625_ (.A(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__o22a_2 _23626_ (.A1(_09180_),
    .A2(_09186_),
    .B1(_09179_),
    .B2(_09187_),
    .X(_09290_));
 sky130_vsdinv _23627_ (.A(_09290_),
    .Y(_09291_));
 sky130_fd_sc_hd__a22o_2 _23628_ (.A1(_09289_),
    .A2(_09290_),
    .B1(_09288_),
    .B2(_09291_),
    .X(_09292_));
 sky130_fd_sc_hd__a2bb2o_2 _23629_ (.A1_N(_09271_),
    .A2_N(_09292_),
    .B1(_09271_),
    .B2(_09292_),
    .X(_09293_));
 sky130_fd_sc_hd__a2bb2o_2 _23630_ (.A1_N(_09274_),
    .A2_N(_09293_),
    .B1(_09274_),
    .B2(_09293_),
    .X(_09294_));
 sky130_fd_sc_hd__a2bb2o_2 _23631_ (.A1_N(_09273_),
    .A2_N(_09294_),
    .B1(_09273_),
    .B2(_09294_),
    .X(_09295_));
 sky130_fd_sc_hd__o22a_2 _23632_ (.A1(_09205_),
    .A2(_09206_),
    .B1(_09200_),
    .B2(_09207_),
    .X(_09296_));
 sky130_fd_sc_hd__o22a_2 _23633_ (.A1(_09212_),
    .A2(_09217_),
    .B1(_09211_),
    .B2(_09218_),
    .X(_09297_));
 sky130_fd_sc_hd__buf_1 _23634_ (.A(_08559_),
    .X(_09298_));
 sky130_fd_sc_hd__o22a_2 _23635_ (.A1(_09298_),
    .A2(_07008_),
    .B1(_05660_),
    .B2(_06891_),
    .X(_09299_));
 sky130_fd_sc_hd__and4_2 _23636_ (.A(_11594_),
    .B(_06876_),
    .C(_11599_),
    .D(_11880_),
    .X(_09300_));
 sky130_fd_sc_hd__nor2_2 _23637_ (.A(_09299_),
    .B(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__buf_1 _23638_ (.A(_07285_),
    .X(_09302_));
 sky130_fd_sc_hd__nor2_2 _23639_ (.A(_05563_),
    .B(_09302_),
    .Y(_09303_));
 sky130_fd_sc_hd__a2bb2o_2 _23640_ (.A1_N(_09301_),
    .A2_N(_09303_),
    .B1(_09301_),
    .B2(_09303_),
    .X(_09304_));
 sky130_fd_sc_hd__buf_1 _23641_ (.A(_09103_),
    .X(_09305_));
 sky130_fd_sc_hd__buf_1 _23642_ (.A(_06031_),
    .X(_09306_));
 sky130_fd_sc_hd__o22a_2 _23643_ (.A1(_09305_),
    .A2(_06378_),
    .B1(_09306_),
    .B2(_06882_),
    .X(_09307_));
 sky130_fd_sc_hd__and4_2 _23644_ (.A(_11587_),
    .B(_11894_),
    .C(_11591_),
    .D(_11890_),
    .X(_09308_));
 sky130_fd_sc_hd__nor2_2 _23645_ (.A(_09307_),
    .B(_09308_),
    .Y(_09309_));
 sky130_fd_sc_hd__buf_1 _23646_ (.A(_05927_),
    .X(_09310_));
 sky130_fd_sc_hd__buf_1 _23647_ (.A(_07015_),
    .X(_09311_));
 sky130_fd_sc_hd__nor2_2 _23648_ (.A(_09310_),
    .B(_09311_),
    .Y(_09312_));
 sky130_fd_sc_hd__a2bb2o_2 _23649_ (.A1_N(_09309_),
    .A2_N(_09312_),
    .B1(_09309_),
    .B2(_09312_),
    .X(_09313_));
 sky130_fd_sc_hd__a21oi_2 _23650_ (.A1(_09203_),
    .A2(_09204_),
    .B1(_09202_),
    .Y(_09314_));
 sky130_fd_sc_hd__a2bb2o_2 _23651_ (.A1_N(_09313_),
    .A2_N(_09314_),
    .B1(_09313_),
    .B2(_09314_),
    .X(_09315_));
 sky130_fd_sc_hd__a2bb2o_2 _23652_ (.A1_N(_09304_),
    .A2_N(_09315_),
    .B1(_09304_),
    .B2(_09315_),
    .X(_09316_));
 sky130_fd_sc_hd__a2bb2o_2 _23653_ (.A1_N(_09297_),
    .A2_N(_09316_),
    .B1(_09297_),
    .B2(_09316_),
    .X(_09317_));
 sky130_fd_sc_hd__a2bb2o_2 _23654_ (.A1_N(_09296_),
    .A2_N(_09317_),
    .B1(_09296_),
    .B2(_09317_),
    .X(_09318_));
 sky130_fd_sc_hd__and4_2 _23655_ (.A(_09128_),
    .B(_05429_),
    .C(_11561_),
    .D(_11913_),
    .X(_09319_));
 sky130_fd_sc_hd__buf_1 _23656_ (.A(_07247_),
    .X(_09320_));
 sky130_fd_sc_hd__o22a_2 _23657_ (.A1(_10597_),
    .A2(_11915_),
    .B1(_09320_),
    .B2(_05510_),
    .X(_09321_));
 sky130_fd_sc_hd__nor2_2 _23658_ (.A(_09319_),
    .B(_09321_),
    .Y(_09322_));
 sky130_fd_sc_hd__nor2_2 _23659_ (.A(_07101_),
    .B(_05704_),
    .Y(_09323_));
 sky130_fd_sc_hd__a2bb2o_2 _23660_ (.A1_N(_09322_),
    .A2_N(_09323_),
    .B1(_09322_),
    .B2(_09323_),
    .X(_09324_));
 sky130_fd_sc_hd__a21oi_2 _23661_ (.A1(_09222_),
    .A2(_09223_),
    .B1(_09220_),
    .Y(_09325_));
 sky130_fd_sc_hd__o2bb2ai_2 _23662_ (.A1_N(_09324_),
    .A2_N(_09325_),
    .B1(_09324_),
    .B2(_09325_),
    .Y(_09326_));
 sky130_fd_sc_hd__o22a_2 _23663_ (.A1(_08917_),
    .A2(_05816_),
    .B1(_06830_),
    .B2(_05885_),
    .X(_09327_));
 sky130_fd_sc_hd__and4_2 _23664_ (.A(_11567_),
    .B(_11909_),
    .C(_11572_),
    .D(_11906_),
    .X(_09328_));
 sky130_fd_sc_hd__nor2_2 _23665_ (.A(_09327_),
    .B(_09328_),
    .Y(_09329_));
 sky130_fd_sc_hd__buf_1 _23666_ (.A(_06687_),
    .X(_09330_));
 sky130_fd_sc_hd__nor2_2 _23667_ (.A(_09330_),
    .B(_05988_),
    .Y(_09331_));
 sky130_fd_sc_hd__a2bb2o_2 _23668_ (.A1_N(_09329_),
    .A2_N(_09331_),
    .B1(_09329_),
    .B2(_09331_),
    .X(_09332_));
 sky130_fd_sc_hd__o2bb2ai_2 _23669_ (.A1_N(_09326_),
    .A2_N(_09332_),
    .B1(_09326_),
    .B2(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__o22a_2 _23670_ (.A1(_09224_),
    .A2(_09225_),
    .B1(_09227_),
    .B2(_09232_),
    .X(_09334_));
 sky130_fd_sc_hd__o2bb2a_2 _23671_ (.A1_N(_09333_),
    .A2_N(_09334_),
    .B1(_09333_),
    .B2(_09334_),
    .X(_09335_));
 sky130_vsdinv _23672_ (.A(_09335_),
    .Y(_09336_));
 sky130_fd_sc_hd__a21oi_2 _23673_ (.A1(_09215_),
    .A2(_09216_),
    .B1(_09214_),
    .Y(_09337_));
 sky130_fd_sc_hd__a21oi_2 _23674_ (.A1(_09230_),
    .A2(_09231_),
    .B1(_09229_),
    .Y(_09338_));
 sky130_fd_sc_hd__buf_1 _23675_ (.A(_08909_),
    .X(_09339_));
 sky130_fd_sc_hd__o22a_2 _23676_ (.A1(_09339_),
    .A2(_06103_),
    .B1(_06443_),
    .B2(_06226_),
    .X(_09340_));
 sky130_fd_sc_hd__and4_2 _23677_ (.A(_11577_),
    .B(_11901_),
    .C(_11582_),
    .D(_11898_),
    .X(_09341_));
 sky130_fd_sc_hd__nor2_2 _23678_ (.A(_09340_),
    .B(_09341_),
    .Y(_09342_));
 sky130_fd_sc_hd__nor2_2 _23679_ (.A(_06275_),
    .B(_06620_),
    .Y(_09343_));
 sky130_fd_sc_hd__a2bb2o_2 _23680_ (.A1_N(_09342_),
    .A2_N(_09343_),
    .B1(_09342_),
    .B2(_09343_),
    .X(_09344_));
 sky130_fd_sc_hd__a2bb2o_2 _23681_ (.A1_N(_09338_),
    .A2_N(_09344_),
    .B1(_09338_),
    .B2(_09344_),
    .X(_09345_));
 sky130_fd_sc_hd__a2bb2o_2 _23682_ (.A1_N(_09337_),
    .A2_N(_09345_),
    .B1(_09337_),
    .B2(_09345_),
    .X(_09346_));
 sky130_vsdinv _23683_ (.A(_09346_),
    .Y(_09347_));
 sky130_fd_sc_hd__a22o_2 _23684_ (.A1(_09336_),
    .A2(_09346_),
    .B1(_09335_),
    .B2(_09347_),
    .X(_09348_));
 sky130_fd_sc_hd__o22a_2 _23685_ (.A1(_09234_),
    .A2(_09235_),
    .B1(_09219_),
    .B2(_09236_),
    .X(_09349_));
 sky130_fd_sc_hd__a2bb2o_2 _23686_ (.A1_N(_09348_),
    .A2_N(_09349_),
    .B1(_09348_),
    .B2(_09349_),
    .X(_09350_));
 sky130_fd_sc_hd__a2bb2o_2 _23687_ (.A1_N(_09318_),
    .A2_N(_09350_),
    .B1(_09318_),
    .B2(_09350_),
    .X(_09351_));
 sky130_fd_sc_hd__o22a_2 _23688_ (.A1(_09237_),
    .A2(_09238_),
    .B1(_09210_),
    .B2(_09239_),
    .X(_09352_));
 sky130_fd_sc_hd__a2bb2o_2 _23689_ (.A1_N(_09351_),
    .A2_N(_09352_),
    .B1(_09351_),
    .B2(_09352_),
    .X(_09353_));
 sky130_fd_sc_hd__a2bb2o_2 _23690_ (.A1_N(_09295_),
    .A2_N(_09353_),
    .B1(_09295_),
    .B2(_09353_),
    .X(_09354_));
 sky130_fd_sc_hd__o22a_2 _23691_ (.A1(_09240_),
    .A2(_09241_),
    .B1(_09193_),
    .B2(_09242_),
    .X(_09355_));
 sky130_fd_sc_hd__a2bb2o_2 _23692_ (.A1_N(_09354_),
    .A2_N(_09355_),
    .B1(_09354_),
    .B2(_09355_),
    .X(_09356_));
 sky130_fd_sc_hd__a2bb2o_2 _23693_ (.A1_N(_09270_),
    .A2_N(_09356_),
    .B1(_09270_),
    .B2(_09356_),
    .X(_09357_));
 sky130_fd_sc_hd__o22a_2 _23694_ (.A1(_09243_),
    .A2(_09244_),
    .B1(_09174_),
    .B2(_09245_),
    .X(_09358_));
 sky130_fd_sc_hd__a2bb2o_2 _23695_ (.A1_N(_09357_),
    .A2_N(_09358_),
    .B1(_09357_),
    .B2(_09358_),
    .X(_09359_));
 sky130_fd_sc_hd__a2bb2o_2 _23696_ (.A1_N(_09261_),
    .A2_N(_09359_),
    .B1(_09261_),
    .B2(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__o22a_2 _23697_ (.A1(_09246_),
    .A2(_09247_),
    .B1(_09163_),
    .B2(_09248_),
    .X(_09361_));
 sky130_fd_sc_hd__a2bb2o_2 _23698_ (.A1_N(_09360_),
    .A2_N(_09361_),
    .B1(_09360_),
    .B2(_09361_),
    .X(_09362_));
 sky130_fd_sc_hd__a2bb2o_2 _23699_ (.A1_N(_09162_),
    .A2_N(_09362_),
    .B1(_09162_),
    .B2(_09362_),
    .X(_09363_));
 sky130_fd_sc_hd__o22a_2 _23700_ (.A1(_09249_),
    .A2(_09250_),
    .B1(_09061_),
    .B2(_09251_),
    .X(_09364_));
 sky130_fd_sc_hd__or2_2 _23701_ (.A(_09363_),
    .B(_09364_),
    .X(_09365_));
 sky130_fd_sc_hd__a21bo_2 _23702_ (.A1(_09363_),
    .A2(_09364_),
    .B1_N(_09365_),
    .X(_09366_));
 sky130_fd_sc_hd__or2_2 _23703_ (.A(_09157_),
    .B(_09255_),
    .X(_09367_));
 sky130_fd_sc_hd__or3_2 _23704_ (.A(_08951_),
    .B(_09058_),
    .C(_09367_),
    .X(_09368_));
 sky130_fd_sc_hd__or2_2 _23705_ (.A(_08953_),
    .B(_09368_),
    .X(_09369_));
 sky130_fd_sc_hd__o221a_2 _23706_ (.A1(_09156_),
    .A2(_09253_),
    .B1(_09158_),
    .B2(_09367_),
    .C1(_09254_),
    .X(_09370_));
 sky130_fd_sc_hd__o221a_2 _23707_ (.A1(_08954_),
    .A2(_09368_),
    .B1(_08502_),
    .B2(_09369_),
    .C1(_09370_),
    .X(_09371_));
 sky130_fd_sc_hd__o31a_2 _23708_ (.A1(_08499_),
    .A2(_09369_),
    .A3(_07425_),
    .B1(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__a2bb2oi_2 _23709_ (.A1_N(_09366_),
    .A2_N(_09372_),
    .B1(_09366_),
    .B2(_09372_),
    .Y(_02667_));
 sky130_fd_sc_hd__o21ai_2 _23710_ (.A1(_09366_),
    .A2(_09372_),
    .B1(_09365_),
    .Y(_09373_));
 sky130_fd_sc_hd__o22a_2 _23711_ (.A1(_09264_),
    .A2(_09268_),
    .B1(_09263_),
    .B2(_09269_),
    .X(_09374_));
 sky130_fd_sc_hd__or2_2 _23712_ (.A(_08842_),
    .B(_09374_),
    .X(_09375_));
 sky130_fd_sc_hd__a21bo_2 _23713_ (.A1(_09258_),
    .A2(_09374_),
    .B1_N(_09375_),
    .X(_09376_));
 sky130_fd_sc_hd__or3_2 _23714_ (.A(_08743_),
    .B(_08850_),
    .C(_09265_),
    .X(_09377_));
 sky130_fd_sc_hd__o21a_2 _23715_ (.A1(_09262_),
    .A2(_09267_),
    .B1(_09377_),
    .X(_09378_));
 sky130_fd_sc_hd__o22a_2 _23716_ (.A1(_09274_),
    .A2(_09293_),
    .B1(_09273_),
    .B2(_09294_),
    .X(_09379_));
 sky130_fd_sc_hd__nand2_2 _23717_ (.A(_09168_),
    .B(_09265_),
    .Y(_09380_));
 sky130_vsdinv _23718_ (.A(_08378_),
    .Y(_09381_));
 sky130_fd_sc_hd__nand2_2 _23719_ (.A(_09377_),
    .B(_09380_),
    .Y(_09382_));
 sky130_fd_sc_hd__a32o_2 _23720_ (.A1(_09377_),
    .A2(_09380_),
    .A3(_09381_),
    .B1(_08623_),
    .B2(_09382_),
    .X(_09383_));
 sky130_fd_sc_hd__buf_1 _23721_ (.A(_09383_),
    .X(_09384_));
 sky130_fd_sc_hd__a2bb2o_2 _23722_ (.A1_N(_09379_),
    .A2_N(_09384_),
    .B1(_09379_),
    .B2(_09384_),
    .X(_09385_));
 sky130_fd_sc_hd__a2bb2o_2 _23723_ (.A1_N(_09378_),
    .A2_N(_09385_),
    .B1(_09378_),
    .B2(_09385_),
    .X(_09386_));
 sky130_fd_sc_hd__o22a_2 _23724_ (.A1(_09289_),
    .A2(_09290_),
    .B1(_09272_),
    .B2(_09292_),
    .X(_09387_));
 sky130_fd_sc_hd__o22a_2 _23725_ (.A1(_09297_),
    .A2(_09316_),
    .B1(_09296_),
    .B2(_09317_),
    .X(_09388_));
 sky130_fd_sc_hd__buf_1 _23726_ (.A(_09178_),
    .X(_09389_));
 sky130_fd_sc_hd__a21oi_2 _23727_ (.A1(_09301_),
    .A2(_09303_),
    .B1(_09300_),
    .Y(_09390_));
 sky130_fd_sc_hd__or4_2 _23728_ (.A(_07727_),
    .B(_06549_),
    .C(_07727_),
    .D(_06428_),
    .X(_09391_));
 sky130_fd_sc_hd__o22a_2 _23729_ (.A1(_10586_),
    .A2(_05389_),
    .B1(_10586_),
    .B2(_07918_),
    .X(_09392_));
 sky130_vsdinv _23730_ (.A(_09392_),
    .Y(_09393_));
 sky130_vsdinv _23731_ (.A(_09391_),
    .Y(_09394_));
 sky130_fd_sc_hd__or2_2 _23732_ (.A(_09394_),
    .B(_09392_),
    .X(_09395_));
 sky130_fd_sc_hd__a32o_2 _23733_ (.A1(_09391_),
    .A2(_09393_),
    .A3(_09185_),
    .B1(_09184_),
    .B2(_09395_),
    .X(_09396_));
 sky130_fd_sc_hd__o2bb2a_2 _23734_ (.A1_N(_09390_),
    .A2_N(_09396_),
    .B1(_09390_),
    .B2(_09396_),
    .X(_09397_));
 sky130_fd_sc_hd__a31o_2 _23735_ (.A1(_09284_),
    .A2(\pcpi_mul.rs2[15] ),
    .A3(_09279_),
    .B1(_09277_),
    .X(_09398_));
 sky130_vsdinv _23736_ (.A(_09397_),
    .Y(_09399_));
 sky130_vsdinv _23737_ (.A(_09398_),
    .Y(_09400_));
 sky130_fd_sc_hd__o22a_2 _23738_ (.A1(_09397_),
    .A2(_09398_),
    .B1(_09399_),
    .B2(_09400_),
    .X(_09401_));
 sky130_vsdinv _23739_ (.A(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__o22a_2 _23740_ (.A1(_09281_),
    .A2(_09282_),
    .B1(_09286_),
    .B2(_09287_),
    .X(_09403_));
 sky130_vsdinv _23741_ (.A(_09403_),
    .Y(_09404_));
 sky130_fd_sc_hd__a22o_2 _23742_ (.A1(_09402_),
    .A2(_09403_),
    .B1(_09401_),
    .B2(_09404_),
    .X(_09405_));
 sky130_fd_sc_hd__a2bb2o_2 _23743_ (.A1_N(_09389_),
    .A2_N(_09405_),
    .B1(_09271_),
    .B2(_09405_),
    .X(_09406_));
 sky130_fd_sc_hd__a2bb2o_2 _23744_ (.A1_N(_09388_),
    .A2_N(_09406_),
    .B1(_09388_),
    .B2(_09406_),
    .X(_09407_));
 sky130_fd_sc_hd__a2bb2o_2 _23745_ (.A1_N(_09387_),
    .A2_N(_09407_),
    .B1(_09387_),
    .B2(_09407_),
    .X(_09408_));
 sky130_fd_sc_hd__and4_2 _23746_ (.A(_09128_),
    .B(_05598_),
    .C(_11561_),
    .D(_05999_),
    .X(_09409_));
 sky130_fd_sc_hd__o22a_2 _23747_ (.A1(_10597_),
    .A2(_11913_),
    .B1(_09320_),
    .B2(_06255_),
    .X(_09410_));
 sky130_fd_sc_hd__nor2_2 _23748_ (.A(_09409_),
    .B(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__nor2_2 _23749_ (.A(_07101_),
    .B(_05816_),
    .Y(_09412_));
 sky130_fd_sc_hd__a2bb2o_2 _23750_ (.A1_N(_09411_),
    .A2_N(_09412_),
    .B1(_09411_),
    .B2(_09412_),
    .X(_09413_));
 sky130_fd_sc_hd__a21oi_2 _23751_ (.A1(_09322_),
    .A2(_09323_),
    .B1(_09319_),
    .Y(_09414_));
 sky130_fd_sc_hd__o2bb2ai_2 _23752_ (.A1_N(_09413_),
    .A2_N(_09414_),
    .B1(_09413_),
    .B2(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__o22a_2 _23753_ (.A1(_08917_),
    .A2(_05824_),
    .B1(_06830_),
    .B2(_05893_),
    .X(_09416_));
 sky130_fd_sc_hd__and4_2 _23754_ (.A(_11567_),
    .B(_11906_),
    .C(_11571_),
    .D(_11903_),
    .X(_09417_));
 sky130_fd_sc_hd__nor2_2 _23755_ (.A(_09416_),
    .B(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__nor2_2 _23756_ (.A(_06687_),
    .B(_06103_),
    .Y(_09419_));
 sky130_fd_sc_hd__a2bb2o_2 _23757_ (.A1_N(_09418_),
    .A2_N(_09419_),
    .B1(_09418_),
    .B2(_09419_),
    .X(_09420_));
 sky130_fd_sc_hd__o2bb2ai_2 _23758_ (.A1_N(_09415_),
    .A2_N(_09420_),
    .B1(_09415_),
    .B2(_09420_),
    .Y(_09421_));
 sky130_fd_sc_hd__o22a_2 _23759_ (.A1(_09324_),
    .A2(_09325_),
    .B1(_09326_),
    .B2(_09332_),
    .X(_09422_));
 sky130_fd_sc_hd__o2bb2ai_2 _23760_ (.A1_N(_09421_),
    .A2_N(_09422_),
    .B1(_09421_),
    .B2(_09422_),
    .Y(_09423_));
 sky130_fd_sc_hd__a21oi_2 _23761_ (.A1(_09342_),
    .A2(_09343_),
    .B1(_09341_),
    .Y(_09424_));
 sky130_fd_sc_hd__a21oi_2 _23762_ (.A1(_09329_),
    .A2(_09331_),
    .B1(_09328_),
    .Y(_09425_));
 sky130_fd_sc_hd__o22a_2 _23763_ (.A1(_09339_),
    .A2(_06360_),
    .B1(_06446_),
    .B2(_06362_),
    .X(_09426_));
 sky130_fd_sc_hd__and4_2 _23764_ (.A(_11576_),
    .B(_11898_),
    .C(_11581_),
    .D(_11896_),
    .X(_09427_));
 sky130_fd_sc_hd__nor2_2 _23765_ (.A(_09426_),
    .B(_09427_),
    .Y(_09428_));
 sky130_fd_sc_hd__buf_1 _23766_ (.A(_06617_),
    .X(_09429_));
 sky130_fd_sc_hd__nor2_2 _23767_ (.A(_06274_),
    .B(_09429_),
    .Y(_09430_));
 sky130_fd_sc_hd__a2bb2o_2 _23768_ (.A1_N(_09428_),
    .A2_N(_09430_),
    .B1(_09428_),
    .B2(_09430_),
    .X(_09431_));
 sky130_fd_sc_hd__a2bb2o_2 _23769_ (.A1_N(_09425_),
    .A2_N(_09431_),
    .B1(_09425_),
    .B2(_09431_),
    .X(_09432_));
 sky130_fd_sc_hd__a2bb2o_2 _23770_ (.A1_N(_09424_),
    .A2_N(_09432_),
    .B1(_09424_),
    .B2(_09432_),
    .X(_09433_));
 sky130_fd_sc_hd__o2bb2ai_2 _23771_ (.A1_N(_09423_),
    .A2_N(_09433_),
    .B1(_09423_),
    .B2(_09433_),
    .Y(_09434_));
 sky130_fd_sc_hd__o22a_2 _23772_ (.A1(_09333_),
    .A2(_09334_),
    .B1(_09336_),
    .B2(_09346_),
    .X(_09435_));
 sky130_fd_sc_hd__o2bb2a_2 _23773_ (.A1_N(_09434_),
    .A2_N(_09435_),
    .B1(_09434_),
    .B2(_09435_),
    .X(_09436_));
 sky130_vsdinv _23774_ (.A(_09436_),
    .Y(_09437_));
 sky130_fd_sc_hd__o22a_2 _23775_ (.A1(_09313_),
    .A2(_09314_),
    .B1(_09304_),
    .B2(_09315_),
    .X(_09438_));
 sky130_fd_sc_hd__o22a_2 _23776_ (.A1(_09338_),
    .A2(_09344_),
    .B1(_09337_),
    .B2(_09345_),
    .X(_09439_));
 sky130_fd_sc_hd__o22a_2 _23777_ (.A1(_09298_),
    .A2(_07010_),
    .B1(_05660_),
    .B2(_07024_),
    .X(_09440_));
 sky130_fd_sc_hd__and4_2 _23778_ (.A(_11594_),
    .B(_07012_),
    .C(_11599_),
    .D(_11878_),
    .X(_09441_));
 sky130_fd_sc_hd__nor2_2 _23779_ (.A(_09440_),
    .B(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__nor2_2 _23780_ (.A(_05563_),
    .B(_07583_),
    .Y(_09443_));
 sky130_fd_sc_hd__a2bb2o_2 _23781_ (.A1_N(_09442_),
    .A2_N(_09443_),
    .B1(_09442_),
    .B2(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__o22a_2 _23782_ (.A1(_09305_),
    .A2(_06882_),
    .B1(_09306_),
    .B2(_07015_),
    .X(_09445_));
 sky130_fd_sc_hd__and4_2 _23783_ (.A(_11587_),
    .B(_11889_),
    .C(_11591_),
    .D(_11886_),
    .X(_09446_));
 sky130_fd_sc_hd__nor2_2 _23784_ (.A(_09445_),
    .B(_09446_),
    .Y(_09447_));
 sky130_fd_sc_hd__nor2_2 _23785_ (.A(_09310_),
    .B(_07151_),
    .Y(_09448_));
 sky130_fd_sc_hd__a2bb2o_2 _23786_ (.A1_N(_09447_),
    .A2_N(_09448_),
    .B1(_09447_),
    .B2(_09448_),
    .X(_09449_));
 sky130_fd_sc_hd__a21oi_2 _23787_ (.A1(_09309_),
    .A2(_09312_),
    .B1(_09308_),
    .Y(_09450_));
 sky130_fd_sc_hd__a2bb2o_2 _23788_ (.A1_N(_09449_),
    .A2_N(_09450_),
    .B1(_09449_),
    .B2(_09450_),
    .X(_09451_));
 sky130_fd_sc_hd__a2bb2o_2 _23789_ (.A1_N(_09444_),
    .A2_N(_09451_),
    .B1(_09444_),
    .B2(_09451_),
    .X(_09452_));
 sky130_fd_sc_hd__a2bb2o_2 _23790_ (.A1_N(_09439_),
    .A2_N(_09452_),
    .B1(_09439_),
    .B2(_09452_),
    .X(_09453_));
 sky130_fd_sc_hd__a2bb2o_2 _23791_ (.A1_N(_09438_),
    .A2_N(_09453_),
    .B1(_09438_),
    .B2(_09453_),
    .X(_09454_));
 sky130_vsdinv _23792_ (.A(_09454_),
    .Y(_09455_));
 sky130_fd_sc_hd__a22o_2 _23793_ (.A1(_09437_),
    .A2(_09454_),
    .B1(_09436_),
    .B2(_09455_),
    .X(_09456_));
 sky130_fd_sc_hd__o22a_2 _23794_ (.A1(_09348_),
    .A2(_09349_),
    .B1(_09318_),
    .B2(_09350_),
    .X(_09457_));
 sky130_fd_sc_hd__a2bb2o_2 _23795_ (.A1_N(_09456_),
    .A2_N(_09457_),
    .B1(_09456_),
    .B2(_09457_),
    .X(_09458_));
 sky130_fd_sc_hd__a2bb2o_2 _23796_ (.A1_N(_09408_),
    .A2_N(_09458_),
    .B1(_09408_),
    .B2(_09458_),
    .X(_09459_));
 sky130_fd_sc_hd__o22a_2 _23797_ (.A1(_09351_),
    .A2(_09352_),
    .B1(_09295_),
    .B2(_09353_),
    .X(_09460_));
 sky130_fd_sc_hd__a2bb2o_2 _23798_ (.A1_N(_09459_),
    .A2_N(_09460_),
    .B1(_09459_),
    .B2(_09460_),
    .X(_09461_));
 sky130_fd_sc_hd__a2bb2o_2 _23799_ (.A1_N(_09386_),
    .A2_N(_09461_),
    .B1(_09386_),
    .B2(_09461_),
    .X(_09462_));
 sky130_fd_sc_hd__o22a_2 _23800_ (.A1(_09354_),
    .A2(_09355_),
    .B1(_09270_),
    .B2(_09356_),
    .X(_09463_));
 sky130_fd_sc_hd__a2bb2o_2 _23801_ (.A1_N(_09462_),
    .A2_N(_09463_),
    .B1(_09462_),
    .B2(_09463_),
    .X(_09464_));
 sky130_fd_sc_hd__a2bb2o_2 _23802_ (.A1_N(_09376_),
    .A2_N(_09464_),
    .B1(_09376_),
    .B2(_09464_),
    .X(_09465_));
 sky130_fd_sc_hd__o22a_2 _23803_ (.A1(_09357_),
    .A2(_09358_),
    .B1(_09261_),
    .B2(_09359_),
    .X(_09466_));
 sky130_fd_sc_hd__a2bb2o_2 _23804_ (.A1_N(_09465_),
    .A2_N(_09466_),
    .B1(_09465_),
    .B2(_09466_),
    .X(_09467_));
 sky130_fd_sc_hd__a2bb2o_2 _23805_ (.A1_N(_09260_),
    .A2_N(_09467_),
    .B1(_09260_),
    .B2(_09467_),
    .X(_09468_));
 sky130_fd_sc_hd__o22a_2 _23806_ (.A1(_09360_),
    .A2(_09361_),
    .B1(_09162_),
    .B2(_09362_),
    .X(_09469_));
 sky130_fd_sc_hd__or2_2 _23807_ (.A(_09468_),
    .B(_09469_),
    .X(_09470_));
 sky130_fd_sc_hd__a21bo_2 _23808_ (.A1(_09468_),
    .A2(_09469_),
    .B1_N(_09470_),
    .X(_09471_));
 sky130_fd_sc_hd__a2bb2o_2 _23809_ (.A1_N(_09373_),
    .A2_N(_09471_),
    .B1(_09373_),
    .B2(_09471_),
    .X(_02668_));
 sky130_fd_sc_hd__buf_1 _23810_ (.A(_09384_),
    .X(_09472_));
 sky130_fd_sc_hd__o22a_2 _23811_ (.A1(_09379_),
    .A2(_09472_),
    .B1(_09378_),
    .B2(_09385_),
    .X(_09473_));
 sky130_fd_sc_hd__or2_2 _23812_ (.A(_08842_),
    .B(_09473_),
    .X(_09474_));
 sky130_fd_sc_hd__a21bo_2 _23813_ (.A1(_09258_),
    .A2(_09473_),
    .B1_N(_09474_),
    .X(_09475_));
 sky130_fd_sc_hd__o21a_2 _23814_ (.A1(_09262_),
    .A2(_09382_),
    .B1(_09377_),
    .X(_09476_));
 sky130_fd_sc_hd__buf_1 _23815_ (.A(_09476_),
    .X(_09477_));
 sky130_fd_sc_hd__buf_1 _23816_ (.A(_09383_),
    .X(_09478_));
 sky130_fd_sc_hd__o22a_2 _23817_ (.A1(_09388_),
    .A2(_09406_),
    .B1(_09387_),
    .B2(_09407_),
    .X(_09479_));
 sky130_fd_sc_hd__a2bb2o_2 _23818_ (.A1_N(_09478_),
    .A2_N(_09479_),
    .B1(_09478_),
    .B2(_09479_),
    .X(_09480_));
 sky130_fd_sc_hd__a2bb2o_2 _23819_ (.A1_N(_09477_),
    .A2_N(_09480_),
    .B1(_09477_),
    .B2(_09480_),
    .X(_09481_));
 sky130_fd_sc_hd__and4_2 _23820_ (.A(_09128_),
    .B(_05607_),
    .C(_11561_),
    .D(_11909_),
    .X(_09482_));
 sky130_fd_sc_hd__o22a_2 _23821_ (.A1(_10597_),
    .A2(_11911_),
    .B1(_09320_),
    .B2(_05716_),
    .X(_09483_));
 sky130_fd_sc_hd__nor2_2 _23822_ (.A(_09482_),
    .B(_09483_),
    .Y(_09484_));
 sky130_fd_sc_hd__nor2_2 _23823_ (.A(_07101_),
    .B(_05885_),
    .Y(_09485_));
 sky130_fd_sc_hd__a2bb2o_2 _23824_ (.A1_N(_09484_),
    .A2_N(_09485_),
    .B1(_09484_),
    .B2(_09485_),
    .X(_09486_));
 sky130_fd_sc_hd__a21oi_2 _23825_ (.A1(_09411_),
    .A2(_09412_),
    .B1(_09409_),
    .Y(_09487_));
 sky130_fd_sc_hd__o2bb2ai_2 _23826_ (.A1_N(_09486_),
    .A2_N(_09487_),
    .B1(_09486_),
    .B2(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__o22a_2 _23827_ (.A1(_08917_),
    .A2(_05893_),
    .B1(_06830_),
    .B2(_08057_),
    .X(_09489_));
 sky130_fd_sc_hd__and4_2 _23828_ (.A(_11567_),
    .B(_11903_),
    .C(_11571_),
    .D(_11900_),
    .X(_09490_));
 sky130_fd_sc_hd__nor2_2 _23829_ (.A(_09489_),
    .B(_09490_),
    .Y(_09491_));
 sky130_fd_sc_hd__nor2_2 _23830_ (.A(_09330_),
    .B(_06226_),
    .Y(_09492_));
 sky130_fd_sc_hd__a2bb2o_2 _23831_ (.A1_N(_09491_),
    .A2_N(_09492_),
    .B1(_09491_),
    .B2(_09492_),
    .X(_09493_));
 sky130_fd_sc_hd__o2bb2ai_2 _23832_ (.A1_N(_09488_),
    .A2_N(_09493_),
    .B1(_09488_),
    .B2(_09493_),
    .Y(_09494_));
 sky130_fd_sc_hd__o22a_2 _23833_ (.A1(_09413_),
    .A2(_09414_),
    .B1(_09415_),
    .B2(_09420_),
    .X(_09495_));
 sky130_fd_sc_hd__o2bb2ai_2 _23834_ (.A1_N(_09494_),
    .A2_N(_09495_),
    .B1(_09494_),
    .B2(_09495_),
    .Y(_09496_));
 sky130_fd_sc_hd__a21oi_2 _23835_ (.A1(_09428_),
    .A2(_09430_),
    .B1(_09427_),
    .Y(_09497_));
 sky130_fd_sc_hd__a21oi_2 _23836_ (.A1(_09418_),
    .A2(_09419_),
    .B1(_09417_),
    .Y(_09498_));
 sky130_fd_sc_hd__o22a_2 _23837_ (.A1(_09339_),
    .A2(_06234_),
    .B1(_06446_),
    .B2(_06617_),
    .X(_09499_));
 sky130_fd_sc_hd__and4_2 _23838_ (.A(_11576_),
    .B(_11895_),
    .C(_11581_),
    .D(_11893_),
    .X(_09500_));
 sky130_fd_sc_hd__nor2_2 _23839_ (.A(_09499_),
    .B(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__nor2_2 _23840_ (.A(_06274_),
    .B(_06882_),
    .Y(_09502_));
 sky130_fd_sc_hd__a2bb2o_2 _23841_ (.A1_N(_09501_),
    .A2_N(_09502_),
    .B1(_09501_),
    .B2(_09502_),
    .X(_09503_));
 sky130_fd_sc_hd__a2bb2o_2 _23842_ (.A1_N(_09498_),
    .A2_N(_09503_),
    .B1(_09498_),
    .B2(_09503_),
    .X(_09504_));
 sky130_fd_sc_hd__a2bb2o_2 _23843_ (.A1_N(_09497_),
    .A2_N(_09504_),
    .B1(_09497_),
    .B2(_09504_),
    .X(_09505_));
 sky130_fd_sc_hd__o2bb2ai_2 _23844_ (.A1_N(_09496_),
    .A2_N(_09505_),
    .B1(_09496_),
    .B2(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__o22a_2 _23845_ (.A1(_09421_),
    .A2(_09422_),
    .B1(_09423_),
    .B2(_09433_),
    .X(_09507_));
 sky130_fd_sc_hd__o2bb2a_2 _23846_ (.A1_N(_09506_),
    .A2_N(_09507_),
    .B1(_09506_),
    .B2(_09507_),
    .X(_09508_));
 sky130_vsdinv _23847_ (.A(_09508_),
    .Y(_09509_));
 sky130_fd_sc_hd__o22a_2 _23848_ (.A1(_09449_),
    .A2(_09450_),
    .B1(_09444_),
    .B2(_09451_),
    .X(_09510_));
 sky130_fd_sc_hd__o22a_2 _23849_ (.A1(_09425_),
    .A2(_09431_),
    .B1(_09424_),
    .B2(_09432_),
    .X(_09511_));
 sky130_fd_sc_hd__o22a_2 _23850_ (.A1(_09298_),
    .A2(_07024_),
    .B1(_05660_),
    .B2(_07160_),
    .X(_09512_));
 sky130_fd_sc_hd__and4_2 _23851_ (.A(_11594_),
    .B(_11878_),
    .C(_11599_),
    .D(_11874_),
    .X(_09513_));
 sky130_fd_sc_hd__or2_2 _23852_ (.A(_09512_),
    .B(_09513_),
    .X(_09514_));
 sky130_vsdinv _23853_ (.A(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__or2_2 _23854_ (.A(_07728_),
    .B(_08437_),
    .X(_09516_));
 sky130_fd_sc_hd__buf_1 _23855_ (.A(_09516_),
    .X(_09517_));
 sky130_fd_sc_hd__a32o_2 _23856_ (.A1(_09284_),
    .A2(\pcpi_mul.rs2[18] ),
    .A3(_09515_),
    .B1(_09514_),
    .B2(_09517_),
    .X(_09518_));
 sky130_fd_sc_hd__o22a_2 _23857_ (.A1(_09305_),
    .A2(_07015_),
    .B1(_09306_),
    .B2(_07151_),
    .X(_09519_));
 sky130_fd_sc_hd__and4_2 _23858_ (.A(_11587_),
    .B(_11885_),
    .C(_11591_),
    .D(_06876_),
    .X(_09520_));
 sky130_fd_sc_hd__nor2_2 _23859_ (.A(_09519_),
    .B(_09520_),
    .Y(_09521_));
 sky130_fd_sc_hd__nor2_2 _23860_ (.A(_09310_),
    .B(_07289_),
    .Y(_09522_));
 sky130_fd_sc_hd__a2bb2o_2 _23861_ (.A1_N(_09521_),
    .A2_N(_09522_),
    .B1(_09521_),
    .B2(_09522_),
    .X(_09523_));
 sky130_fd_sc_hd__a21oi_2 _23862_ (.A1(_09447_),
    .A2(_09448_),
    .B1(_09446_),
    .Y(_09524_));
 sky130_fd_sc_hd__a2bb2o_2 _23863_ (.A1_N(_09523_),
    .A2_N(_09524_),
    .B1(_09523_),
    .B2(_09524_),
    .X(_09525_));
 sky130_fd_sc_hd__a2bb2o_2 _23864_ (.A1_N(_09518_),
    .A2_N(_09525_),
    .B1(_09518_),
    .B2(_09525_),
    .X(_09526_));
 sky130_fd_sc_hd__a2bb2o_2 _23865_ (.A1_N(_09511_),
    .A2_N(_09526_),
    .B1(_09511_),
    .B2(_09526_),
    .X(_09527_));
 sky130_fd_sc_hd__a2bb2o_2 _23866_ (.A1_N(_09510_),
    .A2_N(_09527_),
    .B1(_09510_),
    .B2(_09527_),
    .X(_09528_));
 sky130_vsdinv _23867_ (.A(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__a22o_2 _23868_ (.A1(_09509_),
    .A2(_09528_),
    .B1(_09508_),
    .B2(_09529_),
    .X(_09530_));
 sky130_fd_sc_hd__o22a_2 _23869_ (.A1(_09434_),
    .A2(_09435_),
    .B1(_09437_),
    .B2(_09454_),
    .X(_09531_));
 sky130_fd_sc_hd__a2bb2o_2 _23870_ (.A1_N(_09530_),
    .A2_N(_09531_),
    .B1(_09530_),
    .B2(_09531_),
    .X(_09532_));
 sky130_fd_sc_hd__o22a_2 _23871_ (.A1(_09402_),
    .A2(_09403_),
    .B1(_09272_),
    .B2(_09405_),
    .X(_09533_));
 sky130_fd_sc_hd__o22a_2 _23872_ (.A1(_09439_),
    .A2(_09452_),
    .B1(_09438_),
    .B2(_09453_),
    .X(_09534_));
 sky130_fd_sc_hd__a21oi_2 _23873_ (.A1(_09442_),
    .A2(_09443_),
    .B1(_09441_),
    .Y(_09535_));
 sky130_fd_sc_hd__a2bb2o_2 _23874_ (.A1_N(_09396_),
    .A2_N(_09535_),
    .B1(_09396_),
    .B2(_09535_),
    .X(_09536_));
 sky130_fd_sc_hd__o21a_2 _23875_ (.A1(_09184_),
    .A2(_09395_),
    .B1(_09391_),
    .X(_09537_));
 sky130_fd_sc_hd__buf_1 _23876_ (.A(_09537_),
    .X(_09538_));
 sky130_fd_sc_hd__o2bb2a_2 _23877_ (.A1_N(_09536_),
    .A2_N(_09538_),
    .B1(_09536_),
    .B2(_09538_),
    .X(_09539_));
 sky130_vsdinv _23878_ (.A(_09539_),
    .Y(_09540_));
 sky130_fd_sc_hd__buf_1 _23879_ (.A(_09396_),
    .X(_09541_));
 sky130_fd_sc_hd__o22a_2 _23880_ (.A1(_09390_),
    .A2(_09541_),
    .B1(_09399_),
    .B2(_09400_),
    .X(_09542_));
 sky130_vsdinv _23881_ (.A(_09542_),
    .Y(_09543_));
 sky130_fd_sc_hd__a22o_2 _23882_ (.A1(_09540_),
    .A2(_09542_),
    .B1(_09539_),
    .B2(_09543_),
    .X(_09544_));
 sky130_fd_sc_hd__a2bb2o_2 _23883_ (.A1_N(_09389_),
    .A2_N(_09544_),
    .B1(_09389_),
    .B2(_09544_),
    .X(_09545_));
 sky130_fd_sc_hd__a2bb2o_2 _23884_ (.A1_N(_09534_),
    .A2_N(_09545_),
    .B1(_09534_),
    .B2(_09545_),
    .X(_09546_));
 sky130_fd_sc_hd__a2bb2o_2 _23885_ (.A1_N(_09533_),
    .A2_N(_09546_),
    .B1(_09533_),
    .B2(_09546_),
    .X(_09547_));
 sky130_fd_sc_hd__a2bb2o_2 _23886_ (.A1_N(_09532_),
    .A2_N(_09547_),
    .B1(_09532_),
    .B2(_09547_),
    .X(_09548_));
 sky130_fd_sc_hd__o22a_2 _23887_ (.A1(_09456_),
    .A2(_09457_),
    .B1(_09408_),
    .B2(_09458_),
    .X(_09549_));
 sky130_fd_sc_hd__a2bb2o_2 _23888_ (.A1_N(_09548_),
    .A2_N(_09549_),
    .B1(_09548_),
    .B2(_09549_),
    .X(_09550_));
 sky130_fd_sc_hd__a2bb2o_2 _23889_ (.A1_N(_09481_),
    .A2_N(_09550_),
    .B1(_09481_),
    .B2(_09550_),
    .X(_09551_));
 sky130_fd_sc_hd__o22a_2 _23890_ (.A1(_09459_),
    .A2(_09460_),
    .B1(_09386_),
    .B2(_09461_),
    .X(_09552_));
 sky130_fd_sc_hd__a2bb2o_2 _23891_ (.A1_N(_09551_),
    .A2_N(_09552_),
    .B1(_09551_),
    .B2(_09552_),
    .X(_09553_));
 sky130_fd_sc_hd__a2bb2o_2 _23892_ (.A1_N(_09475_),
    .A2_N(_09553_),
    .B1(_09475_),
    .B2(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__o22a_2 _23893_ (.A1(_09462_),
    .A2(_09463_),
    .B1(_09376_),
    .B2(_09464_),
    .X(_09555_));
 sky130_fd_sc_hd__a2bb2o_2 _23894_ (.A1_N(_09554_),
    .A2_N(_09555_),
    .B1(_09554_),
    .B2(_09555_),
    .X(_09556_));
 sky130_fd_sc_hd__a2bb2o_2 _23895_ (.A1_N(_09375_),
    .A2_N(_09556_),
    .B1(_09375_),
    .B2(_09556_),
    .X(_09557_));
 sky130_fd_sc_hd__o22a_2 _23896_ (.A1(_09465_),
    .A2(_09466_),
    .B1(_09260_),
    .B2(_09467_),
    .X(_09558_));
 sky130_fd_sc_hd__or2_2 _23897_ (.A(_09557_),
    .B(_09558_),
    .X(_09559_));
 sky130_fd_sc_hd__a21bo_2 _23898_ (.A1(_09557_),
    .A2(_09558_),
    .B1_N(_09559_),
    .X(_09560_));
 sky130_fd_sc_hd__a22o_2 _23899_ (.A1(_09468_),
    .A2(_09469_),
    .B1(_09365_),
    .B2(_09470_),
    .X(_09561_));
 sky130_fd_sc_hd__o31a_2 _23900_ (.A1(_09366_),
    .A2(_09471_),
    .A3(_09372_),
    .B1(_09561_),
    .X(_09562_));
 sky130_fd_sc_hd__a2bb2oi_2 _23901_ (.A1_N(_09560_),
    .A2_N(_09562_),
    .B1(_09560_),
    .B2(_09562_),
    .Y(_02669_));
 sky130_fd_sc_hd__buf_1 _23902_ (.A(_09384_),
    .X(_09563_));
 sky130_fd_sc_hd__buf_1 _23903_ (.A(_09476_),
    .X(_09564_));
 sky130_fd_sc_hd__o22a_2 _23904_ (.A1(_09563_),
    .A2(_09479_),
    .B1(_09564_),
    .B2(_09480_),
    .X(_09565_));
 sky130_fd_sc_hd__or2_2 _23905_ (.A(_09257_),
    .B(_09565_),
    .X(_09566_));
 sky130_fd_sc_hd__a21bo_2 _23906_ (.A1(_09258_),
    .A2(_09565_),
    .B1_N(_09566_),
    .X(_09567_));
 sky130_fd_sc_hd__and4_2 _23907_ (.A(_09128_),
    .B(_05815_),
    .C(_11561_),
    .D(_06240_),
    .X(_09568_));
 sky130_fd_sc_hd__o22a_2 _23908_ (.A1(_10597_),
    .A2(_11909_),
    .B1(_09320_),
    .B2(_05824_),
    .X(_09569_));
 sky130_fd_sc_hd__nor2_2 _23909_ (.A(_09568_),
    .B(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__nor2_2 _23910_ (.A(_07101_),
    .B(_05988_),
    .Y(_09571_));
 sky130_fd_sc_hd__a2bb2o_2 _23911_ (.A1_N(_09570_),
    .A2_N(_09571_),
    .B1(_09570_),
    .B2(_09571_),
    .X(_09572_));
 sky130_fd_sc_hd__a21oi_2 _23912_ (.A1(_09484_),
    .A2(_09485_),
    .B1(_09482_),
    .Y(_09573_));
 sky130_fd_sc_hd__o2bb2ai_2 _23913_ (.A1_N(_09572_),
    .A2_N(_09573_),
    .B1(_09572_),
    .B2(_09573_),
    .Y(_09574_));
 sky130_fd_sc_hd__o22a_2 _23914_ (.A1(_08917_),
    .A2(_08057_),
    .B1(_06831_),
    .B2(_06360_),
    .X(_09575_));
 sky130_fd_sc_hd__and4_2 _23915_ (.A(_11568_),
    .B(_11901_),
    .C(_11572_),
    .D(_11897_),
    .X(_09576_));
 sky130_fd_sc_hd__nor2_2 _23916_ (.A(_09575_),
    .B(_09576_),
    .Y(_09577_));
 sky130_fd_sc_hd__nor2_2 _23917_ (.A(_09330_),
    .B(_06620_),
    .Y(_09578_));
 sky130_fd_sc_hd__a2bb2o_2 _23918_ (.A1_N(_09577_),
    .A2_N(_09578_),
    .B1(_09577_),
    .B2(_09578_),
    .X(_09579_));
 sky130_fd_sc_hd__o2bb2ai_2 _23919_ (.A1_N(_09574_),
    .A2_N(_09579_),
    .B1(_09574_),
    .B2(_09579_),
    .Y(_09580_));
 sky130_fd_sc_hd__o22a_2 _23920_ (.A1(_09486_),
    .A2(_09487_),
    .B1(_09488_),
    .B2(_09493_),
    .X(_09581_));
 sky130_fd_sc_hd__o2bb2ai_2 _23921_ (.A1_N(_09580_),
    .A2_N(_09581_),
    .B1(_09580_),
    .B2(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__a21oi_2 _23922_ (.A1(_09501_),
    .A2(_09502_),
    .B1(_09500_),
    .Y(_09583_));
 sky130_fd_sc_hd__a21oi_2 _23923_ (.A1(_09491_),
    .A2(_09492_),
    .B1(_09490_),
    .Y(_09584_));
 sky130_fd_sc_hd__o22a_2 _23924_ (.A1(_09339_),
    .A2(_06617_),
    .B1(_06446_),
    .B2(_06497_),
    .X(_09585_));
 sky130_fd_sc_hd__and4_2 _23925_ (.A(_11576_),
    .B(_11893_),
    .C(_11581_),
    .D(_11889_),
    .X(_09586_));
 sky130_fd_sc_hd__nor2_2 _23926_ (.A(_09585_),
    .B(_09586_),
    .Y(_09587_));
 sky130_fd_sc_hd__nor2_2 _23927_ (.A(_06274_),
    .B(_07015_),
    .Y(_09588_));
 sky130_fd_sc_hd__a2bb2o_2 _23928_ (.A1_N(_09587_),
    .A2_N(_09588_),
    .B1(_09587_),
    .B2(_09588_),
    .X(_09589_));
 sky130_fd_sc_hd__a2bb2o_2 _23929_ (.A1_N(_09584_),
    .A2_N(_09589_),
    .B1(_09584_),
    .B2(_09589_),
    .X(_09590_));
 sky130_fd_sc_hd__a2bb2o_2 _23930_ (.A1_N(_09583_),
    .A2_N(_09590_),
    .B1(_09583_),
    .B2(_09590_),
    .X(_09591_));
 sky130_fd_sc_hd__o2bb2ai_2 _23931_ (.A1_N(_09582_),
    .A2_N(_09591_),
    .B1(_09582_),
    .B2(_09591_),
    .Y(_09592_));
 sky130_fd_sc_hd__o22a_2 _23932_ (.A1(_09494_),
    .A2(_09495_),
    .B1(_09496_),
    .B2(_09505_),
    .X(_09593_));
 sky130_fd_sc_hd__o2bb2a_2 _23933_ (.A1_N(_09592_),
    .A2_N(_09593_),
    .B1(_09592_),
    .B2(_09593_),
    .X(_09594_));
 sky130_vsdinv _23934_ (.A(_09594_),
    .Y(_09595_));
 sky130_fd_sc_hd__o22a_2 _23935_ (.A1(_09523_),
    .A2(_09524_),
    .B1(_09518_),
    .B2(_09525_),
    .X(_09596_));
 sky130_fd_sc_hd__o22a_2 _23936_ (.A1(_09498_),
    .A2(_09503_),
    .B1(_09497_),
    .B2(_09504_),
    .X(_09597_));
 sky130_fd_sc_hd__nor2_2 _23937_ (.A(_09298_),
    .B(_07583_),
    .Y(_09598_));
 sky130_fd_sc_hd__or2_2 _23938_ (.A(_10586_),
    .B(_05660_),
    .X(_09599_));
 sky130_vsdinv _23939_ (.A(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__a2bb2o_2 _23940_ (.A1_N(_09598_),
    .A2_N(_09600_),
    .B1(_09598_),
    .B2(_09600_),
    .X(_09601_));
 sky130_fd_sc_hd__a2bb2o_2 _23941_ (.A1_N(_09517_),
    .A2_N(_09601_),
    .B1(_09517_),
    .B2(_09601_),
    .X(_09602_));
 sky130_fd_sc_hd__o22a_2 _23942_ (.A1(_09305_),
    .A2(_07008_),
    .B1(_09306_),
    .B2(_07010_),
    .X(_09603_));
 sky130_fd_sc_hd__and4_2 _23943_ (.A(_11587_),
    .B(_06876_),
    .C(_11591_),
    .D(_07012_),
    .X(_09604_));
 sky130_fd_sc_hd__nor2_2 _23944_ (.A(_09603_),
    .B(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__nor2_2 _23945_ (.A(_05927_),
    .B(_09302_),
    .Y(_09606_));
 sky130_fd_sc_hd__a2bb2o_2 _23946_ (.A1_N(_09605_),
    .A2_N(_09606_),
    .B1(_09605_),
    .B2(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__a21oi_2 _23947_ (.A1(_09521_),
    .A2(_09522_),
    .B1(_09520_),
    .Y(_09608_));
 sky130_fd_sc_hd__a2bb2o_2 _23948_ (.A1_N(_09607_),
    .A2_N(_09608_),
    .B1(_09607_),
    .B2(_09608_),
    .X(_09609_));
 sky130_fd_sc_hd__a2bb2o_2 _23949_ (.A1_N(_09602_),
    .A2_N(_09609_),
    .B1(_09602_),
    .B2(_09609_),
    .X(_09610_));
 sky130_fd_sc_hd__a2bb2o_2 _23950_ (.A1_N(_09597_),
    .A2_N(_09610_),
    .B1(_09597_),
    .B2(_09610_),
    .X(_09611_));
 sky130_fd_sc_hd__a2bb2o_2 _23951_ (.A1_N(_09596_),
    .A2_N(_09611_),
    .B1(_09596_),
    .B2(_09611_),
    .X(_09612_));
 sky130_vsdinv _23952_ (.A(_09612_),
    .Y(_09613_));
 sky130_fd_sc_hd__a22o_2 _23953_ (.A1(_09595_),
    .A2(_09612_),
    .B1(_09594_),
    .B2(_09613_),
    .X(_09614_));
 sky130_fd_sc_hd__o22a_2 _23954_ (.A1(_09506_),
    .A2(_09507_),
    .B1(_09509_),
    .B2(_09528_),
    .X(_09615_));
 sky130_fd_sc_hd__a2bb2o_2 _23955_ (.A1_N(_09614_),
    .A2_N(_09615_),
    .B1(_09614_),
    .B2(_09615_),
    .X(_09616_));
 sky130_fd_sc_hd__o22a_2 _23956_ (.A1(_09540_),
    .A2(_09542_),
    .B1(_09272_),
    .B2(_09544_),
    .X(_09617_));
 sky130_fd_sc_hd__o22a_2 _23957_ (.A1(_09511_),
    .A2(_09526_),
    .B1(_09510_),
    .B2(_09527_),
    .X(_09618_));
 sky130_fd_sc_hd__o21ba_2 _23958_ (.A1(_09514_),
    .A2(_09517_),
    .B1_N(_09513_),
    .X(_09619_));
 sky130_fd_sc_hd__a2bb2o_2 _23959_ (.A1_N(_09541_),
    .A2_N(_09619_),
    .B1(_09541_),
    .B2(_09619_),
    .X(_09620_));
 sky130_fd_sc_hd__a2bb2o_2 _23960_ (.A1_N(_09538_),
    .A2_N(_09620_),
    .B1(_09538_),
    .B2(_09620_),
    .X(_09621_));
 sky130_fd_sc_hd__o22a_2 _23961_ (.A1(_09541_),
    .A2(_09535_),
    .B1(_09536_),
    .B2(_09538_),
    .X(_09622_));
 sky130_fd_sc_hd__o2bb2ai_2 _23962_ (.A1_N(_09621_),
    .A2_N(_09622_),
    .B1(_09621_),
    .B2(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__a2bb2o_2 _23963_ (.A1_N(_09271_),
    .A2_N(_09623_),
    .B1(_09271_),
    .B2(_09623_),
    .X(_09624_));
 sky130_fd_sc_hd__a2bb2o_2 _23964_ (.A1_N(_09618_),
    .A2_N(_09624_),
    .B1(_09618_),
    .B2(_09624_),
    .X(_09625_));
 sky130_fd_sc_hd__a2bb2o_2 _23965_ (.A1_N(_09617_),
    .A2_N(_09625_),
    .B1(_09617_),
    .B2(_09625_),
    .X(_09626_));
 sky130_fd_sc_hd__a2bb2o_2 _23966_ (.A1_N(_09616_),
    .A2_N(_09626_),
    .B1(_09616_),
    .B2(_09626_),
    .X(_09627_));
 sky130_fd_sc_hd__o22a_2 _23967_ (.A1(_09530_),
    .A2(_09531_),
    .B1(_09532_),
    .B2(_09547_),
    .X(_09628_));
 sky130_fd_sc_hd__a2bb2o_2 _23968_ (.A1_N(_09627_),
    .A2_N(_09628_),
    .B1(_09627_),
    .B2(_09628_),
    .X(_09629_));
 sky130_fd_sc_hd__buf_1 _23969_ (.A(_09476_),
    .X(_09630_));
 sky130_fd_sc_hd__o22a_2 _23970_ (.A1(_09534_),
    .A2(_09545_),
    .B1(_09533_),
    .B2(_09546_),
    .X(_09631_));
 sky130_fd_sc_hd__a2bb2o_2 _23971_ (.A1_N(_09472_),
    .A2_N(_09631_),
    .B1(_09472_),
    .B2(_09631_),
    .X(_09632_));
 sky130_fd_sc_hd__a2bb2o_2 _23972_ (.A1_N(_09630_),
    .A2_N(_09632_),
    .B1(_09630_),
    .B2(_09632_),
    .X(_09633_));
 sky130_fd_sc_hd__a2bb2o_2 _23973_ (.A1_N(_09629_),
    .A2_N(_09633_),
    .B1(_09629_),
    .B2(_09633_),
    .X(_09634_));
 sky130_fd_sc_hd__o22a_2 _23974_ (.A1(_09548_),
    .A2(_09549_),
    .B1(_09481_),
    .B2(_09550_),
    .X(_09635_));
 sky130_fd_sc_hd__a2bb2o_2 _23975_ (.A1_N(_09634_),
    .A2_N(_09635_),
    .B1(_09634_),
    .B2(_09635_),
    .X(_09636_));
 sky130_fd_sc_hd__a2bb2o_2 _23976_ (.A1_N(_09567_),
    .A2_N(_09636_),
    .B1(_09567_),
    .B2(_09636_),
    .X(_09637_));
 sky130_fd_sc_hd__o22a_2 _23977_ (.A1(_09551_),
    .A2(_09552_),
    .B1(_09475_),
    .B2(_09553_),
    .X(_09638_));
 sky130_fd_sc_hd__a2bb2o_2 _23978_ (.A1_N(_09637_),
    .A2_N(_09638_),
    .B1(_09637_),
    .B2(_09638_),
    .X(_09639_));
 sky130_fd_sc_hd__a2bb2o_2 _23979_ (.A1_N(_09474_),
    .A2_N(_09639_),
    .B1(_09474_),
    .B2(_09639_),
    .X(_09640_));
 sky130_fd_sc_hd__o22a_2 _23980_ (.A1(_09554_),
    .A2(_09555_),
    .B1(_09375_),
    .B2(_09556_),
    .X(_09641_));
 sky130_fd_sc_hd__and2_2 _23981_ (.A(_09640_),
    .B(_09641_),
    .X(_09642_));
 sky130_fd_sc_hd__or2_2 _23982_ (.A(_09640_),
    .B(_09641_),
    .X(_09643_));
 sky130_fd_sc_hd__or2b_2 _23983_ (.A(_09642_),
    .B_N(_09643_),
    .X(_09644_));
 sky130_fd_sc_hd__o21ai_2 _23984_ (.A1(_09560_),
    .A2(_09562_),
    .B1(_09559_),
    .Y(_09645_));
 sky130_fd_sc_hd__a2bb2o_2 _23985_ (.A1_N(_09644_),
    .A2_N(_09645_),
    .B1(_09644_),
    .B2(_09645_),
    .X(_02670_));
 sky130_fd_sc_hd__buf_1 _23986_ (.A(_09128_),
    .X(_09646_));
 sky130_fd_sc_hd__and4_2 _23987_ (.A(_09646_),
    .B(_05824_),
    .C(_11561_),
    .D(_06372_),
    .X(_09647_));
 sky130_fd_sc_hd__o22a_2 _23988_ (.A1(_10598_),
    .A2(_11906_),
    .B1(_09320_),
    .B2(_05893_),
    .X(_09648_));
 sky130_fd_sc_hd__nor2_2 _23989_ (.A(_09647_),
    .B(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__buf_1 _23990_ (.A(_07101_),
    .X(_09650_));
 sky130_fd_sc_hd__nor2_2 _23991_ (.A(_09650_),
    .B(_06103_),
    .Y(_09651_));
 sky130_fd_sc_hd__a2bb2o_2 _23992_ (.A1_N(_09649_),
    .A2_N(_09651_),
    .B1(_09649_),
    .B2(_09651_),
    .X(_09652_));
 sky130_fd_sc_hd__a21oi_2 _23993_ (.A1(_09570_),
    .A2(_09571_),
    .B1(_09568_),
    .Y(_09653_));
 sky130_fd_sc_hd__o2bb2ai_2 _23994_ (.A1_N(_09652_),
    .A2_N(_09653_),
    .B1(_09652_),
    .B2(_09653_),
    .Y(_09654_));
 sky130_fd_sc_hd__buf_1 _23995_ (.A(_08917_),
    .X(_09655_));
 sky130_fd_sc_hd__o22a_2 _23996_ (.A1(_09655_),
    .A2(_06226_),
    .B1(_06831_),
    .B2(_06362_),
    .X(_09656_));
 sky130_fd_sc_hd__and4_2 _23997_ (.A(_11568_),
    .B(_11898_),
    .C(_11572_),
    .D(_11896_),
    .X(_09657_));
 sky130_fd_sc_hd__nor2_2 _23998_ (.A(_09656_),
    .B(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__nor2_2 _23999_ (.A(_09330_),
    .B(_09429_),
    .Y(_09659_));
 sky130_fd_sc_hd__a2bb2o_2 _24000_ (.A1_N(_09658_),
    .A2_N(_09659_),
    .B1(_09658_),
    .B2(_09659_),
    .X(_09660_));
 sky130_fd_sc_hd__o2bb2ai_2 _24001_ (.A1_N(_09654_),
    .A2_N(_09660_),
    .B1(_09654_),
    .B2(_09660_),
    .Y(_09661_));
 sky130_fd_sc_hd__o22a_2 _24002_ (.A1(_09572_),
    .A2(_09573_),
    .B1(_09574_),
    .B2(_09579_),
    .X(_09662_));
 sky130_fd_sc_hd__o2bb2ai_2 _24003_ (.A1_N(_09661_),
    .A2_N(_09662_),
    .B1(_09661_),
    .B2(_09662_),
    .Y(_09663_));
 sky130_fd_sc_hd__a21oi_2 _24004_ (.A1(_09587_),
    .A2(_09588_),
    .B1(_09586_),
    .Y(_09664_));
 sky130_fd_sc_hd__a21oi_2 _24005_ (.A1(_09577_),
    .A2(_09578_),
    .B1(_09576_),
    .Y(_09665_));
 sky130_fd_sc_hd__o22a_2 _24006_ (.A1(_09339_),
    .A2(_06882_),
    .B1(_06446_),
    .B2(_06625_),
    .X(_09666_));
 sky130_fd_sc_hd__and4_2 _24007_ (.A(_11576_),
    .B(_11889_),
    .C(_11581_),
    .D(_11885_),
    .X(_09667_));
 sky130_fd_sc_hd__nor2_2 _24008_ (.A(_09666_),
    .B(_09667_),
    .Y(_09668_));
 sky130_fd_sc_hd__nor2_2 _24009_ (.A(_06274_),
    .B(_07151_),
    .Y(_09669_));
 sky130_fd_sc_hd__a2bb2o_2 _24010_ (.A1_N(_09668_),
    .A2_N(_09669_),
    .B1(_09668_),
    .B2(_09669_),
    .X(_09670_));
 sky130_fd_sc_hd__a2bb2o_2 _24011_ (.A1_N(_09665_),
    .A2_N(_09670_),
    .B1(_09665_),
    .B2(_09670_),
    .X(_09671_));
 sky130_fd_sc_hd__a2bb2o_2 _24012_ (.A1_N(_09664_),
    .A2_N(_09671_),
    .B1(_09664_),
    .B2(_09671_),
    .X(_09672_));
 sky130_fd_sc_hd__o2bb2ai_2 _24013_ (.A1_N(_09663_),
    .A2_N(_09672_),
    .B1(_09663_),
    .B2(_09672_),
    .Y(_09673_));
 sky130_fd_sc_hd__o22a_2 _24014_ (.A1(_09580_),
    .A2(_09581_),
    .B1(_09582_),
    .B2(_09591_),
    .X(_09674_));
 sky130_fd_sc_hd__o2bb2ai_2 _24015_ (.A1_N(_09673_),
    .A2_N(_09674_),
    .B1(_09673_),
    .B2(_09674_),
    .Y(_09675_));
 sky130_fd_sc_hd__o22a_2 _24016_ (.A1(_09607_),
    .A2(_09608_),
    .B1(_09602_),
    .B2(_09609_),
    .X(_09676_));
 sky130_fd_sc_hd__o22a_2 _24017_ (.A1(_09584_),
    .A2(_09589_),
    .B1(_09583_),
    .B2(_09590_),
    .X(_09677_));
 sky130_fd_sc_hd__or2_2 _24018_ (.A(_07728_),
    .B(_09298_),
    .X(_09678_));
 sky130_fd_sc_hd__a32o_2 _24019_ (.A1(_07870_),
    .A2(_11594_),
    .A3(_09600_),
    .B1(_09599_),
    .B2(_09678_),
    .X(_09679_));
 sky130_fd_sc_hd__a2bb2o_2 _24020_ (.A1_N(_09516_),
    .A2_N(_09679_),
    .B1(_09516_),
    .B2(_09679_),
    .X(_09680_));
 sky130_fd_sc_hd__o22a_2 _24021_ (.A1(_09103_),
    .A2(_06891_),
    .B1(_06031_),
    .B2(_07285_),
    .X(_09681_));
 sky130_fd_sc_hd__and4_2 _24022_ (.A(_11586_),
    .B(_11880_),
    .C(_11590_),
    .D(_11877_),
    .X(_09682_));
 sky130_fd_sc_hd__nor2_2 _24023_ (.A(_09681_),
    .B(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__nor2_2 _24024_ (.A(_09310_),
    .B(_07583_),
    .Y(_09684_));
 sky130_fd_sc_hd__a2bb2o_2 _24025_ (.A1_N(_09683_),
    .A2_N(_09684_),
    .B1(_09683_),
    .B2(_09684_),
    .X(_09685_));
 sky130_fd_sc_hd__a21oi_2 _24026_ (.A1(_09605_),
    .A2(_09606_),
    .B1(_09604_),
    .Y(_09686_));
 sky130_fd_sc_hd__a2bb2o_2 _24027_ (.A1_N(_09685_),
    .A2_N(_09686_),
    .B1(_09685_),
    .B2(_09686_),
    .X(_09687_));
 sky130_fd_sc_hd__a2bb2o_2 _24028_ (.A1_N(_09680_),
    .A2_N(_09687_),
    .B1(_09680_),
    .B2(_09687_),
    .X(_09688_));
 sky130_fd_sc_hd__a2bb2o_2 _24029_ (.A1_N(_09677_),
    .A2_N(_09688_),
    .B1(_09677_),
    .B2(_09688_),
    .X(_09689_));
 sky130_fd_sc_hd__a2bb2o_2 _24030_ (.A1_N(_09676_),
    .A2_N(_09689_),
    .B1(_09676_),
    .B2(_09689_),
    .X(_09690_));
 sky130_fd_sc_hd__o2bb2ai_2 _24031_ (.A1_N(_09675_),
    .A2_N(_09690_),
    .B1(_09675_),
    .B2(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__o22a_2 _24032_ (.A1(_09592_),
    .A2(_09593_),
    .B1(_09595_),
    .B2(_09612_),
    .X(_09692_));
 sky130_fd_sc_hd__o2bb2a_2 _24033_ (.A1_N(_09691_),
    .A2_N(_09692_),
    .B1(_09691_),
    .B2(_09692_),
    .X(_09693_));
 sky130_vsdinv _24034_ (.A(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__o22a_2 _24035_ (.A1(_09621_),
    .A2(_09622_),
    .B1(_09389_),
    .B2(_09623_),
    .X(_09695_));
 sky130_fd_sc_hd__o22a_2 _24036_ (.A1(_09597_),
    .A2(_09610_),
    .B1(_09596_),
    .B2(_09611_),
    .X(_09696_));
 sky130_fd_sc_hd__buf_1 _24037_ (.A(_09178_),
    .X(_09697_));
 sky130_fd_sc_hd__o22a_2 _24038_ (.A1(_09541_),
    .A2(_09619_),
    .B1(_09538_),
    .B2(_09620_),
    .X(_09698_));
 sky130_fd_sc_hd__buf_1 _24039_ (.A(_07583_),
    .X(_09699_));
 sky130_fd_sc_hd__o32a_2 _24040_ (.A1(_09298_),
    .A2(_09699_),
    .A3(_09599_),
    .B1(_09517_),
    .B2(_09601_),
    .X(_09700_));
 sky130_vsdinv _24041_ (.A(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__nor2_2 _24042_ (.A(_09185_),
    .B(_09393_),
    .Y(_09702_));
 sky130_fd_sc_hd__a21oi_2 _24043_ (.A1(\pcpi_mul.rs2[15] ),
    .A2(_09394_),
    .B1(_09702_),
    .Y(_09703_));
 sky130_fd_sc_hd__a2bb2o_2 _24044_ (.A1_N(_09701_),
    .A2_N(_09703_),
    .B1(_09701_),
    .B2(_09703_),
    .X(_09704_));
 sky130_fd_sc_hd__o2bb2ai_2 _24045_ (.A1_N(_09698_),
    .A2_N(_09704_),
    .B1(_09698_),
    .B2(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__a2bb2o_2 _24046_ (.A1_N(_09697_),
    .A2_N(_09705_),
    .B1(_09697_),
    .B2(_09705_),
    .X(_09706_));
 sky130_fd_sc_hd__a2bb2o_2 _24047_ (.A1_N(_09696_),
    .A2_N(_09706_),
    .B1(_09696_),
    .B2(_09706_),
    .X(_09707_));
 sky130_fd_sc_hd__a2bb2o_2 _24048_ (.A1_N(_09695_),
    .A2_N(_09707_),
    .B1(_09695_),
    .B2(_09707_),
    .X(_09708_));
 sky130_vsdinv _24049_ (.A(_09708_),
    .Y(_09709_));
 sky130_fd_sc_hd__a22o_2 _24050_ (.A1(_09694_),
    .A2(_09708_),
    .B1(_09693_),
    .B2(_09709_),
    .X(_09710_));
 sky130_fd_sc_hd__o22a_2 _24051_ (.A1(_09614_),
    .A2(_09615_),
    .B1(_09616_),
    .B2(_09626_),
    .X(_09711_));
 sky130_fd_sc_hd__a2bb2o_2 _24052_ (.A1_N(_09710_),
    .A2_N(_09711_),
    .B1(_09710_),
    .B2(_09711_),
    .X(_09712_));
 sky130_fd_sc_hd__o22a_2 _24053_ (.A1(_09618_),
    .A2(_09624_),
    .B1(_09617_),
    .B2(_09625_),
    .X(_09713_));
 sky130_fd_sc_hd__a2bb2o_2 _24054_ (.A1_N(_09478_),
    .A2_N(_09713_),
    .B1(_09478_),
    .B2(_09713_),
    .X(_09714_));
 sky130_fd_sc_hd__a2bb2o_2 _24055_ (.A1_N(_09477_),
    .A2_N(_09714_),
    .B1(_09477_),
    .B2(_09714_),
    .X(_09715_));
 sky130_fd_sc_hd__a2bb2o_2 _24056_ (.A1_N(_09712_),
    .A2_N(_09715_),
    .B1(_09712_),
    .B2(_09715_),
    .X(_09716_));
 sky130_fd_sc_hd__o22a_2 _24057_ (.A1(_09627_),
    .A2(_09628_),
    .B1(_09629_),
    .B2(_09633_),
    .X(_09717_));
 sky130_fd_sc_hd__a2bb2o_2 _24058_ (.A1_N(_09716_),
    .A2_N(_09717_),
    .B1(_09716_),
    .B2(_09717_),
    .X(_09718_));
 sky130_fd_sc_hd__buf_1 _24059_ (.A(_09257_),
    .X(_09719_));
 sky130_fd_sc_hd__o22a_2 _24060_ (.A1(_09563_),
    .A2(_09631_),
    .B1(_09564_),
    .B2(_09632_),
    .X(_09720_));
 sky130_fd_sc_hd__or2_2 _24061_ (.A(_09257_),
    .B(_09720_),
    .X(_09721_));
 sky130_fd_sc_hd__a21bo_2 _24062_ (.A1(_09719_),
    .A2(_09720_),
    .B1_N(_09721_),
    .X(_09722_));
 sky130_fd_sc_hd__a2bb2o_2 _24063_ (.A1_N(_09718_),
    .A2_N(_09722_),
    .B1(_09718_),
    .B2(_09722_),
    .X(_09723_));
 sky130_fd_sc_hd__o22a_2 _24064_ (.A1(_09634_),
    .A2(_09635_),
    .B1(_09567_),
    .B2(_09636_),
    .X(_09724_));
 sky130_fd_sc_hd__a2bb2o_2 _24065_ (.A1_N(_09723_),
    .A2_N(_09724_),
    .B1(_09723_),
    .B2(_09724_),
    .X(_09725_));
 sky130_fd_sc_hd__a2bb2o_2 _24066_ (.A1_N(_09566_),
    .A2_N(_09725_),
    .B1(_09566_),
    .B2(_09725_),
    .X(_09726_));
 sky130_fd_sc_hd__o22a_2 _24067_ (.A1(_09637_),
    .A2(_09638_),
    .B1(_09474_),
    .B2(_09639_),
    .X(_09727_));
 sky130_fd_sc_hd__or2_2 _24068_ (.A(_09726_),
    .B(_09727_),
    .X(_09728_));
 sky130_fd_sc_hd__a21bo_2 _24069_ (.A1(_09726_),
    .A2(_09727_),
    .B1_N(_09728_),
    .X(_09729_));
 sky130_fd_sc_hd__or2_2 _24070_ (.A(_09560_),
    .B(_09644_),
    .X(_09730_));
 sky130_fd_sc_hd__or3_2 _24071_ (.A(_09366_),
    .B(_09471_),
    .C(_09730_),
    .X(_09731_));
 sky130_fd_sc_hd__o221a_2 _24072_ (.A1(_09559_),
    .A2(_09642_),
    .B1(_09561_),
    .B2(_09730_),
    .C1(_09643_),
    .X(_09732_));
 sky130_fd_sc_hd__o21ai_2 _24073_ (.A1(_09372_),
    .A2(_09731_),
    .B1(_09732_),
    .Y(_09733_));
 sky130_vsdinv _24074_ (.A(_09733_),
    .Y(_09734_));
 sky130_vsdinv _24075_ (.A(_09729_),
    .Y(_09735_));
 sky130_fd_sc_hd__o22a_2 _24076_ (.A1(_09729_),
    .A2(_09734_),
    .B1(_09735_),
    .B2(_09733_),
    .X(_02671_));
 sky130_fd_sc_hd__o21ai_2 _24077_ (.A1(_09729_),
    .A2(_09734_),
    .B1(_09728_),
    .Y(_09736_));
 sky130_fd_sc_hd__and4_2 _24078_ (.A(_09646_),
    .B(_05987_),
    .C(_11562_),
    .D(_11900_),
    .X(_09737_));
 sky130_fd_sc_hd__buf_1 _24079_ (.A(_09320_),
    .X(_09738_));
 sky130_fd_sc_hd__o22a_2 _24080_ (.A1(_10598_),
    .A2(_11903_),
    .B1(_09738_),
    .B2(_08057_),
    .X(_09739_));
 sky130_fd_sc_hd__nor2_2 _24081_ (.A(_09737_),
    .B(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__nor2_2 _24082_ (.A(_09650_),
    .B(_06226_),
    .Y(_09741_));
 sky130_fd_sc_hd__a2bb2o_2 _24083_ (.A1_N(_09740_),
    .A2_N(_09741_),
    .B1(_09740_),
    .B2(_09741_),
    .X(_09742_));
 sky130_fd_sc_hd__a21oi_2 _24084_ (.A1(_09649_),
    .A2(_09651_),
    .B1(_09647_),
    .Y(_09743_));
 sky130_fd_sc_hd__o2bb2ai_2 _24085_ (.A1_N(_09742_),
    .A2_N(_09743_),
    .B1(_09742_),
    .B2(_09743_),
    .Y(_09744_));
 sky130_fd_sc_hd__o22a_2 _24086_ (.A1(_09655_),
    .A2(_06620_),
    .B1(_06831_),
    .B2(_06378_),
    .X(_09745_));
 sky130_fd_sc_hd__and4_2 _24087_ (.A(_11568_),
    .B(_11896_),
    .C(_11572_),
    .D(_11894_),
    .X(_09746_));
 sky130_fd_sc_hd__nor2_2 _24088_ (.A(_09745_),
    .B(_09746_),
    .Y(_09747_));
 sky130_fd_sc_hd__buf_1 _24089_ (.A(_06882_),
    .X(_09748_));
 sky130_fd_sc_hd__nor2_2 _24090_ (.A(_09330_),
    .B(_09748_),
    .Y(_09749_));
 sky130_fd_sc_hd__a2bb2o_2 _24091_ (.A1_N(_09747_),
    .A2_N(_09749_),
    .B1(_09747_),
    .B2(_09749_),
    .X(_09750_));
 sky130_fd_sc_hd__o2bb2ai_2 _24092_ (.A1_N(_09744_),
    .A2_N(_09750_),
    .B1(_09744_),
    .B2(_09750_),
    .Y(_09751_));
 sky130_fd_sc_hd__o22a_2 _24093_ (.A1(_09652_),
    .A2(_09653_),
    .B1(_09654_),
    .B2(_09660_),
    .X(_09752_));
 sky130_fd_sc_hd__o2bb2ai_2 _24094_ (.A1_N(_09751_),
    .A2_N(_09752_),
    .B1(_09751_),
    .B2(_09752_),
    .Y(_09753_));
 sky130_fd_sc_hd__a21oi_2 _24095_ (.A1(_09668_),
    .A2(_09669_),
    .B1(_09667_),
    .Y(_09754_));
 sky130_fd_sc_hd__a21oi_2 _24096_ (.A1(_09658_),
    .A2(_09659_),
    .B1(_09657_),
    .Y(_09755_));
 sky130_fd_sc_hd__o22a_2 _24097_ (.A1(_09339_),
    .A2(_06625_),
    .B1(_06446_),
    .B2(_07008_),
    .X(_09756_));
 sky130_fd_sc_hd__and4_2 _24098_ (.A(_11576_),
    .B(_11885_),
    .C(_11582_),
    .D(_06876_),
    .X(_09757_));
 sky130_fd_sc_hd__nor2_2 _24099_ (.A(_09756_),
    .B(_09757_),
    .Y(_09758_));
 sky130_fd_sc_hd__nor2_2 _24100_ (.A(_06274_),
    .B(_07289_),
    .Y(_09759_));
 sky130_fd_sc_hd__a2bb2o_2 _24101_ (.A1_N(_09758_),
    .A2_N(_09759_),
    .B1(_09758_),
    .B2(_09759_),
    .X(_09760_));
 sky130_fd_sc_hd__a2bb2o_2 _24102_ (.A1_N(_09755_),
    .A2_N(_09760_),
    .B1(_09755_),
    .B2(_09760_),
    .X(_09761_));
 sky130_fd_sc_hd__a2bb2o_2 _24103_ (.A1_N(_09754_),
    .A2_N(_09761_),
    .B1(_09754_),
    .B2(_09761_),
    .X(_09762_));
 sky130_fd_sc_hd__o2bb2ai_2 _24104_ (.A1_N(_09753_),
    .A2_N(_09762_),
    .B1(_09753_),
    .B2(_09762_),
    .Y(_09763_));
 sky130_fd_sc_hd__o22a_2 _24105_ (.A1(_09661_),
    .A2(_09662_),
    .B1(_09663_),
    .B2(_09672_),
    .X(_09764_));
 sky130_fd_sc_hd__o2bb2ai_2 _24106_ (.A1_N(_09763_),
    .A2_N(_09764_),
    .B1(_09763_),
    .B2(_09764_),
    .Y(_09765_));
 sky130_fd_sc_hd__buf_1 _24107_ (.A(_09680_),
    .X(_09766_));
 sky130_fd_sc_hd__o22a_2 _24108_ (.A1(_09685_),
    .A2(_09686_),
    .B1(_09766_),
    .B2(_09687_),
    .X(_09767_));
 sky130_fd_sc_hd__o22a_2 _24109_ (.A1(_09665_),
    .A2(_09670_),
    .B1(_09664_),
    .B2(_09671_),
    .X(_09768_));
 sky130_fd_sc_hd__o22a_2 _24110_ (.A1(_09103_),
    .A2(_07285_),
    .B1(_06031_),
    .B2(_08266_),
    .X(_09769_));
 sky130_fd_sc_hd__and4_2 _24111_ (.A(_11586_),
    .B(_11877_),
    .C(_11590_),
    .D(_11874_),
    .X(_09770_));
 sky130_fd_sc_hd__nor2_2 _24112_ (.A(_09769_),
    .B(_09770_),
    .Y(_09771_));
 sky130_fd_sc_hd__or2_2 _24113_ (.A(_07728_),
    .B(_08445_),
    .X(_09772_));
 sky130_vsdinv _24114_ (.A(_09772_),
    .Y(_09773_));
 sky130_fd_sc_hd__a2bb2o_2 _24115_ (.A1_N(_09771_),
    .A2_N(_09773_),
    .B1(_09771_),
    .B2(_09773_),
    .X(_09774_));
 sky130_fd_sc_hd__a31o_2 _24116_ (.A1(\pcpi_mul.rs2[21] ),
    .A2(_11874_),
    .A3(_09683_),
    .B1(_09682_),
    .X(_09775_));
 sky130_vsdinv _24117_ (.A(_09775_),
    .Y(_09776_));
 sky130_vsdinv _24118_ (.A(_09774_),
    .Y(_09777_));
 sky130_fd_sc_hd__a22o_2 _24119_ (.A1(_09774_),
    .A2(_09776_),
    .B1(_09777_),
    .B2(_09775_),
    .X(_09778_));
 sky130_fd_sc_hd__a2bb2o_2 _24120_ (.A1_N(_09680_),
    .A2_N(_09778_),
    .B1(_09680_),
    .B2(_09778_),
    .X(_09779_));
 sky130_fd_sc_hd__a2bb2o_2 _24121_ (.A1_N(_09768_),
    .A2_N(_09779_),
    .B1(_09768_),
    .B2(_09779_),
    .X(_09780_));
 sky130_fd_sc_hd__a2bb2o_2 _24122_ (.A1_N(_09767_),
    .A2_N(_09780_),
    .B1(_09767_),
    .B2(_09780_),
    .X(_09781_));
 sky130_fd_sc_hd__o2bb2ai_2 _24123_ (.A1_N(_09765_),
    .A2_N(_09781_),
    .B1(_09765_),
    .B2(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__o22a_2 _24124_ (.A1(_09673_),
    .A2(_09674_),
    .B1(_09675_),
    .B2(_09690_),
    .X(_09783_));
 sky130_fd_sc_hd__o2bb2a_2 _24125_ (.A1_N(_09782_),
    .A2_N(_09783_),
    .B1(_09782_),
    .B2(_09783_),
    .X(_09784_));
 sky130_vsdinv _24126_ (.A(_09784_),
    .Y(_09785_));
 sky130_fd_sc_hd__o22a_2 _24127_ (.A1(_09698_),
    .A2(_09704_),
    .B1(_09389_),
    .B2(_09705_),
    .X(_09786_));
 sky130_fd_sc_hd__o22a_2 _24128_ (.A1(_09677_),
    .A2(_09688_),
    .B1(_09676_),
    .B2(_09689_),
    .X(_09787_));
 sky130_fd_sc_hd__o22a_2 _24129_ (.A1(_09599_),
    .A2(_09678_),
    .B1(_09517_),
    .B2(_09679_),
    .X(_09788_));
 sky130_fd_sc_hd__o22ai_2 _24130_ (.A1(_05310_),
    .A2(_09391_),
    .B1(_09701_),
    .B2(_09702_),
    .Y(_09789_));
 sky130_fd_sc_hd__o2bb2a_2 _24131_ (.A1_N(_09788_),
    .A2_N(_09789_),
    .B1(_09788_),
    .B2(_09789_),
    .X(_09790_));
 sky130_fd_sc_hd__a2bb2o_2 _24132_ (.A1_N(_09697_),
    .A2_N(_09790_),
    .B1(_09697_),
    .B2(_09790_),
    .X(_09791_));
 sky130_fd_sc_hd__a2bb2o_2 _24133_ (.A1_N(_09787_),
    .A2_N(_09791_),
    .B1(_09787_),
    .B2(_09791_),
    .X(_09792_));
 sky130_fd_sc_hd__a2bb2o_2 _24134_ (.A1_N(_09786_),
    .A2_N(_09792_),
    .B1(_09786_),
    .B2(_09792_),
    .X(_09793_));
 sky130_vsdinv _24135_ (.A(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__a22o_2 _24136_ (.A1(_09785_),
    .A2(_09793_),
    .B1(_09784_),
    .B2(_09794_),
    .X(_09795_));
 sky130_fd_sc_hd__o22a_2 _24137_ (.A1(_09691_),
    .A2(_09692_),
    .B1(_09694_),
    .B2(_09708_),
    .X(_09796_));
 sky130_fd_sc_hd__a2bb2o_2 _24138_ (.A1_N(_09795_),
    .A2_N(_09796_),
    .B1(_09795_),
    .B2(_09796_),
    .X(_09797_));
 sky130_fd_sc_hd__o22a_2 _24139_ (.A1(_09696_),
    .A2(_09706_),
    .B1(_09695_),
    .B2(_09707_),
    .X(_09798_));
 sky130_fd_sc_hd__a2bb2o_2 _24140_ (.A1_N(_09384_),
    .A2_N(_09798_),
    .B1(_09384_),
    .B2(_09798_),
    .X(_09799_));
 sky130_fd_sc_hd__a2bb2o_2 _24141_ (.A1_N(_09477_),
    .A2_N(_09799_),
    .B1(_09477_),
    .B2(_09799_),
    .X(_09800_));
 sky130_fd_sc_hd__a2bb2o_2 _24142_ (.A1_N(_09797_),
    .A2_N(_09800_),
    .B1(_09797_),
    .B2(_09800_),
    .X(_09801_));
 sky130_fd_sc_hd__o22a_2 _24143_ (.A1(_09710_),
    .A2(_09711_),
    .B1(_09712_),
    .B2(_09715_),
    .X(_09802_));
 sky130_fd_sc_hd__a2bb2o_2 _24144_ (.A1_N(_09801_),
    .A2_N(_09802_),
    .B1(_09801_),
    .B2(_09802_),
    .X(_09803_));
 sky130_fd_sc_hd__o22a_2 _24145_ (.A1(_09563_),
    .A2(_09713_),
    .B1(_09564_),
    .B2(_09714_),
    .X(_09804_));
 sky130_fd_sc_hd__or2_2 _24146_ (.A(_08842_),
    .B(_09804_),
    .X(_09805_));
 sky130_fd_sc_hd__a21bo_2 _24147_ (.A1(_09258_),
    .A2(_09804_),
    .B1_N(_09805_),
    .X(_09806_));
 sky130_fd_sc_hd__a2bb2o_2 _24148_ (.A1_N(_09803_),
    .A2_N(_09806_),
    .B1(_09803_),
    .B2(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__o22a_2 _24149_ (.A1(_09716_),
    .A2(_09717_),
    .B1(_09718_),
    .B2(_09722_),
    .X(_09808_));
 sky130_fd_sc_hd__a2bb2o_2 _24150_ (.A1_N(_09807_),
    .A2_N(_09808_),
    .B1(_09807_),
    .B2(_09808_),
    .X(_09809_));
 sky130_fd_sc_hd__a2bb2o_2 _24151_ (.A1_N(_09721_),
    .A2_N(_09809_),
    .B1(_09721_),
    .B2(_09809_),
    .X(_09810_));
 sky130_fd_sc_hd__o22a_2 _24152_ (.A1(_09723_),
    .A2(_09724_),
    .B1(_09566_),
    .B2(_09725_),
    .X(_09811_));
 sky130_fd_sc_hd__or2_2 _24153_ (.A(_09810_),
    .B(_09811_),
    .X(_09812_));
 sky130_fd_sc_hd__a21bo_2 _24154_ (.A1(_09810_),
    .A2(_09811_),
    .B1_N(_09812_),
    .X(_09813_));
 sky130_fd_sc_hd__a2bb2o_2 _24155_ (.A1_N(_09736_),
    .A2_N(_09813_),
    .B1(_09736_),
    .B2(_09813_),
    .X(_02672_));
 sky130_fd_sc_hd__and4_2 _24156_ (.A(_09646_),
    .B(_05996_),
    .C(_11562_),
    .D(_11897_),
    .X(_09814_));
 sky130_fd_sc_hd__o22a_2 _24157_ (.A1(_10598_),
    .A2(_11901_),
    .B1(_09738_),
    .B2(_06360_),
    .X(_09815_));
 sky130_fd_sc_hd__nor2_2 _24158_ (.A(_09814_),
    .B(_09815_),
    .Y(_09816_));
 sky130_fd_sc_hd__nor2_2 _24159_ (.A(_09650_),
    .B(_06620_),
    .Y(_09817_));
 sky130_fd_sc_hd__a2bb2o_2 _24160_ (.A1_N(_09816_),
    .A2_N(_09817_),
    .B1(_09816_),
    .B2(_09817_),
    .X(_09818_));
 sky130_fd_sc_hd__a21oi_2 _24161_ (.A1(_09740_),
    .A2(_09741_),
    .B1(_09737_),
    .Y(_09819_));
 sky130_fd_sc_hd__o2bb2ai_2 _24162_ (.A1_N(_09818_),
    .A2_N(_09819_),
    .B1(_09818_),
    .B2(_09819_),
    .Y(_09820_));
 sky130_fd_sc_hd__o22a_2 _24163_ (.A1(_09655_),
    .A2(_09429_),
    .B1(_06831_),
    .B2(_09748_),
    .X(_09821_));
 sky130_fd_sc_hd__and4_2 _24164_ (.A(_11568_),
    .B(_11894_),
    .C(_11572_),
    .D(_11890_),
    .X(_09822_));
 sky130_fd_sc_hd__nor2_2 _24165_ (.A(_09821_),
    .B(_09822_),
    .Y(_09823_));
 sky130_fd_sc_hd__buf_1 _24166_ (.A(_09330_),
    .X(_09824_));
 sky130_fd_sc_hd__nor2_2 _24167_ (.A(_09824_),
    .B(_09311_),
    .Y(_09825_));
 sky130_fd_sc_hd__a2bb2o_2 _24168_ (.A1_N(_09823_),
    .A2_N(_09825_),
    .B1(_09823_),
    .B2(_09825_),
    .X(_09826_));
 sky130_fd_sc_hd__o2bb2ai_2 _24169_ (.A1_N(_09820_),
    .A2_N(_09826_),
    .B1(_09820_),
    .B2(_09826_),
    .Y(_09827_));
 sky130_fd_sc_hd__o22a_2 _24170_ (.A1(_09742_),
    .A2(_09743_),
    .B1(_09744_),
    .B2(_09750_),
    .X(_09828_));
 sky130_fd_sc_hd__o2bb2ai_2 _24171_ (.A1_N(_09827_),
    .A2_N(_09828_),
    .B1(_09827_),
    .B2(_09828_),
    .Y(_09829_));
 sky130_fd_sc_hd__a21oi_2 _24172_ (.A1(_09758_),
    .A2(_09759_),
    .B1(_09757_),
    .Y(_09830_));
 sky130_fd_sc_hd__a21oi_2 _24173_ (.A1(_09747_),
    .A2(_09749_),
    .B1(_09746_),
    .Y(_09831_));
 sky130_fd_sc_hd__buf_1 _24174_ (.A(_08909_),
    .X(_09832_));
 sky130_fd_sc_hd__o22a_2 _24175_ (.A1(_09832_),
    .A2(_07151_),
    .B1(_06443_),
    .B2(_07010_),
    .X(_09833_));
 sky130_fd_sc_hd__and4_2 _24176_ (.A(_11577_),
    .B(_11883_),
    .C(_11582_),
    .D(_07012_),
    .X(_09834_));
 sky130_fd_sc_hd__nor2_2 _24177_ (.A(_09833_),
    .B(_09834_),
    .Y(_09835_));
 sky130_fd_sc_hd__nor2_2 _24178_ (.A(_06275_),
    .B(_09302_),
    .Y(_09836_));
 sky130_fd_sc_hd__a2bb2o_2 _24179_ (.A1_N(_09835_),
    .A2_N(_09836_),
    .B1(_09835_),
    .B2(_09836_),
    .X(_09837_));
 sky130_fd_sc_hd__a2bb2o_2 _24180_ (.A1_N(_09831_),
    .A2_N(_09837_),
    .B1(_09831_),
    .B2(_09837_),
    .X(_09838_));
 sky130_fd_sc_hd__a2bb2o_2 _24181_ (.A1_N(_09830_),
    .A2_N(_09838_),
    .B1(_09830_),
    .B2(_09838_),
    .X(_09839_));
 sky130_fd_sc_hd__o2bb2ai_2 _24182_ (.A1_N(_09829_),
    .A2_N(_09839_),
    .B1(_09829_),
    .B2(_09839_),
    .Y(_09840_));
 sky130_fd_sc_hd__o22a_2 _24183_ (.A1(_09751_),
    .A2(_09752_),
    .B1(_09753_),
    .B2(_09762_),
    .X(_09841_));
 sky130_fd_sc_hd__o2bb2ai_2 _24184_ (.A1_N(_09840_),
    .A2_N(_09841_),
    .B1(_09840_),
    .B2(_09841_),
    .Y(_09842_));
 sky130_fd_sc_hd__o22a_2 _24185_ (.A1(_09774_),
    .A2(_09776_),
    .B1(_09766_),
    .B2(_09778_),
    .X(_09843_));
 sky130_fd_sc_hd__o22a_2 _24186_ (.A1(_09755_),
    .A2(_09760_),
    .B1(_09754_),
    .B2(_09761_),
    .X(_09844_));
 sky130_fd_sc_hd__a31o_2 _24187_ (.A1(_09284_),
    .A2(\pcpi_mul.rs2[21] ),
    .A3(_09771_),
    .B1(_09770_),
    .X(_09845_));
 sky130_vsdinv _24188_ (.A(_09845_),
    .Y(_09846_));
 sky130_fd_sc_hd__o22a_2 _24189_ (.A1(_09103_),
    .A2(_08266_),
    .B1(_07728_),
    .B2(_06031_),
    .X(_09847_));
 sky130_fd_sc_hd__and4_2 _24190_ (.A(_11587_),
    .B(_11874_),
    .C(_07869_),
    .D(_11591_),
    .X(_09848_));
 sky130_fd_sc_hd__nor2_2 _24191_ (.A(_09847_),
    .B(_09848_),
    .Y(_09849_));
 sky130_fd_sc_hd__o2bb2a_2 _24192_ (.A1_N(_09773_),
    .A2_N(_09849_),
    .B1(_09773_),
    .B2(_09849_),
    .X(_09850_));
 sky130_vsdinv _24193_ (.A(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__a22o_2 _24194_ (.A1(_09846_),
    .A2(_09851_),
    .B1(_09845_),
    .B2(_09850_),
    .X(_09852_));
 sky130_fd_sc_hd__a2bb2o_2 _24195_ (.A1_N(_09766_),
    .A2_N(_09852_),
    .B1(_09680_),
    .B2(_09852_),
    .X(_09853_));
 sky130_fd_sc_hd__a2bb2o_2 _24196_ (.A1_N(_09844_),
    .A2_N(_09853_),
    .B1(_09844_),
    .B2(_09853_),
    .X(_09854_));
 sky130_fd_sc_hd__a2bb2o_2 _24197_ (.A1_N(_09843_),
    .A2_N(_09854_),
    .B1(_09843_),
    .B2(_09854_),
    .X(_09855_));
 sky130_fd_sc_hd__o2bb2ai_2 _24198_ (.A1_N(_09842_),
    .A2_N(_09855_),
    .B1(_09842_),
    .B2(_09855_),
    .Y(_09856_));
 sky130_fd_sc_hd__o22a_2 _24199_ (.A1(_09763_),
    .A2(_09764_),
    .B1(_09765_),
    .B2(_09781_),
    .X(_09857_));
 sky130_fd_sc_hd__o2bb2a_2 _24200_ (.A1_N(_09856_),
    .A2_N(_09857_),
    .B1(_09856_),
    .B2(_09857_),
    .X(_09858_));
 sky130_vsdinv _24201_ (.A(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__or3_2 _24202_ (.A(_05310_),
    .B(_09391_),
    .C(_09788_),
    .X(_09860_));
 sky130_fd_sc_hd__o21a_2 _24203_ (.A1(_09389_),
    .A2(_09790_),
    .B1(_09860_),
    .X(_09861_));
 sky130_fd_sc_hd__o22a_2 _24204_ (.A1(_09768_),
    .A2(_09779_),
    .B1(_09767_),
    .B2(_09780_),
    .X(_09862_));
 sky130_vsdinv _24205_ (.A(_09860_),
    .Y(_09863_));
 sky130_fd_sc_hd__and3_2 _24206_ (.A(_09541_),
    .B(_09788_),
    .C(_09537_),
    .X(_09864_));
 sky130_fd_sc_hd__or2_2 _24207_ (.A(_09863_),
    .B(_09864_),
    .X(_09865_));
 sky130_fd_sc_hd__a2bb2o_2 _24208_ (.A1_N(_09697_),
    .A2_N(_09865_),
    .B1(_09697_),
    .B2(_09865_),
    .X(_09866_));
 sky130_fd_sc_hd__a2bb2o_2 _24209_ (.A1_N(_09862_),
    .A2_N(_09866_),
    .B1(_09862_),
    .B2(_09866_),
    .X(_09867_));
 sky130_fd_sc_hd__a2bb2o_2 _24210_ (.A1_N(_09861_),
    .A2_N(_09867_),
    .B1(_09861_),
    .B2(_09867_),
    .X(_09868_));
 sky130_vsdinv _24211_ (.A(_09868_),
    .Y(_09869_));
 sky130_fd_sc_hd__a22o_2 _24212_ (.A1(_09859_),
    .A2(_09868_),
    .B1(_09858_),
    .B2(_09869_),
    .X(_09870_));
 sky130_fd_sc_hd__o22a_2 _24213_ (.A1(_09782_),
    .A2(_09783_),
    .B1(_09785_),
    .B2(_09793_),
    .X(_09871_));
 sky130_fd_sc_hd__a2bb2o_2 _24214_ (.A1_N(_09870_),
    .A2_N(_09871_),
    .B1(_09870_),
    .B2(_09871_),
    .X(_09872_));
 sky130_fd_sc_hd__o22a_2 _24215_ (.A1(_09787_),
    .A2(_09791_),
    .B1(_09786_),
    .B2(_09792_),
    .X(_09873_));
 sky130_fd_sc_hd__a2bb2o_2 _24216_ (.A1_N(_09478_),
    .A2_N(_09873_),
    .B1(_09478_),
    .B2(_09873_),
    .X(_09874_));
 sky130_fd_sc_hd__a2bb2o_2 _24217_ (.A1_N(_09564_),
    .A2_N(_09874_),
    .B1(_09564_),
    .B2(_09874_),
    .X(_09875_));
 sky130_fd_sc_hd__a2bb2o_2 _24218_ (.A1_N(_09872_),
    .A2_N(_09875_),
    .B1(_09872_),
    .B2(_09875_),
    .X(_09876_));
 sky130_fd_sc_hd__o22a_2 _24219_ (.A1(_09795_),
    .A2(_09796_),
    .B1(_09797_),
    .B2(_09800_),
    .X(_09877_));
 sky130_fd_sc_hd__a2bb2o_2 _24220_ (.A1_N(_09876_),
    .A2_N(_09877_),
    .B1(_09876_),
    .B2(_09877_),
    .X(_09878_));
 sky130_fd_sc_hd__o22a_2 _24221_ (.A1(_09472_),
    .A2(_09798_),
    .B1(_09476_),
    .B2(_09799_),
    .X(_09879_));
 sky130_fd_sc_hd__or2_2 _24222_ (.A(_08842_),
    .B(_09879_),
    .X(_09880_));
 sky130_fd_sc_hd__a21bo_2 _24223_ (.A1(_09258_),
    .A2(_09879_),
    .B1_N(_09880_),
    .X(_09881_));
 sky130_fd_sc_hd__a2bb2o_2 _24224_ (.A1_N(_09878_),
    .A2_N(_09881_),
    .B1(_09878_),
    .B2(_09881_),
    .X(_09882_));
 sky130_fd_sc_hd__o22a_2 _24225_ (.A1(_09801_),
    .A2(_09802_),
    .B1(_09803_),
    .B2(_09806_),
    .X(_09883_));
 sky130_fd_sc_hd__a2bb2o_2 _24226_ (.A1_N(_09882_),
    .A2_N(_09883_),
    .B1(_09882_),
    .B2(_09883_),
    .X(_09884_));
 sky130_fd_sc_hd__a2bb2o_2 _24227_ (.A1_N(_09805_),
    .A2_N(_09884_),
    .B1(_09805_),
    .B2(_09884_),
    .X(_09885_));
 sky130_fd_sc_hd__o22a_2 _24228_ (.A1(_09807_),
    .A2(_09808_),
    .B1(_09721_),
    .B2(_09809_),
    .X(_09886_));
 sky130_fd_sc_hd__or2_2 _24229_ (.A(_09885_),
    .B(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__a21bo_2 _24230_ (.A1(_09885_),
    .A2(_09886_),
    .B1_N(_09887_),
    .X(_09888_));
 sky130_fd_sc_hd__a22o_2 _24231_ (.A1(_09810_),
    .A2(_09811_),
    .B1(_09728_),
    .B2(_09812_),
    .X(_09889_));
 sky130_fd_sc_hd__o31a_2 _24232_ (.A1(_09729_),
    .A2(_09813_),
    .A3(_09734_),
    .B1(_09889_),
    .X(_09890_));
 sky130_fd_sc_hd__a2bb2oi_2 _24233_ (.A1_N(_09888_),
    .A2_N(_09890_),
    .B1(_09888_),
    .B2(_09890_),
    .Y(_02673_));
 sky130_fd_sc_hd__and4_2 _24234_ (.A(_09646_),
    .B(_06360_),
    .C(_11562_),
    .D(_11896_),
    .X(_09891_));
 sky130_fd_sc_hd__o22a_2 _24235_ (.A1(_10598_),
    .A2(_11898_),
    .B1(_09738_),
    .B2(_06362_),
    .X(_09892_));
 sky130_fd_sc_hd__nor2_2 _24236_ (.A(_09891_),
    .B(_09892_),
    .Y(_09893_));
 sky130_fd_sc_hd__nor2_2 _24237_ (.A(_09650_),
    .B(_09429_),
    .Y(_09894_));
 sky130_fd_sc_hd__a2bb2o_2 _24238_ (.A1_N(_09893_),
    .A2_N(_09894_),
    .B1(_09893_),
    .B2(_09894_),
    .X(_09895_));
 sky130_fd_sc_hd__a21oi_2 _24239_ (.A1(_09816_),
    .A2(_09817_),
    .B1(_09814_),
    .Y(_09896_));
 sky130_fd_sc_hd__o2bb2ai_2 _24240_ (.A1_N(_09895_),
    .A2_N(_09896_),
    .B1(_09895_),
    .B2(_09896_),
    .Y(_09897_));
 sky130_fd_sc_hd__buf_1 _24241_ (.A(_06831_),
    .X(_09898_));
 sky130_fd_sc_hd__o22a_2 _24242_ (.A1(_09655_),
    .A2(_09748_),
    .B1(_09898_),
    .B2(_07015_),
    .X(_09899_));
 sky130_fd_sc_hd__and4_2 _24243_ (.A(_11568_),
    .B(_11890_),
    .C(_11573_),
    .D(_11886_),
    .X(_09900_));
 sky130_fd_sc_hd__nor2_2 _24244_ (.A(_09899_),
    .B(_09900_),
    .Y(_09901_));
 sky130_fd_sc_hd__buf_1 _24245_ (.A(_07151_),
    .X(_09902_));
 sky130_fd_sc_hd__nor2_2 _24246_ (.A(_09824_),
    .B(_09902_),
    .Y(_09903_));
 sky130_fd_sc_hd__a2bb2o_2 _24247_ (.A1_N(_09901_),
    .A2_N(_09903_),
    .B1(_09901_),
    .B2(_09903_),
    .X(_09904_));
 sky130_fd_sc_hd__o2bb2ai_2 _24248_ (.A1_N(_09897_),
    .A2_N(_09904_),
    .B1(_09897_),
    .B2(_09904_),
    .Y(_09905_));
 sky130_fd_sc_hd__o22a_2 _24249_ (.A1(_09818_),
    .A2(_09819_),
    .B1(_09820_),
    .B2(_09826_),
    .X(_09906_));
 sky130_fd_sc_hd__o2bb2ai_2 _24250_ (.A1_N(_09905_),
    .A2_N(_09906_),
    .B1(_09905_),
    .B2(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__a21oi_2 _24251_ (.A1(_09835_),
    .A2(_09836_),
    .B1(_09834_),
    .Y(_09908_));
 sky130_fd_sc_hd__a21oi_2 _24252_ (.A1(_09823_),
    .A2(_09825_),
    .B1(_09822_),
    .Y(_09909_));
 sky130_fd_sc_hd__o22a_2 _24253_ (.A1(_09832_),
    .A2(_07289_),
    .B1(_06443_),
    .B2(_09302_),
    .X(_09910_));
 sky130_fd_sc_hd__and4_2 _24254_ (.A(_11577_),
    .B(_11881_),
    .C(_11582_),
    .D(_11878_),
    .X(_09911_));
 sky130_fd_sc_hd__nor2_2 _24255_ (.A(_09910_),
    .B(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__nor2_2 _24256_ (.A(_06275_),
    .B(_09699_),
    .Y(_09913_));
 sky130_fd_sc_hd__a2bb2o_2 _24257_ (.A1_N(_09912_),
    .A2_N(_09913_),
    .B1(_09912_),
    .B2(_09913_),
    .X(_09914_));
 sky130_fd_sc_hd__a2bb2o_2 _24258_ (.A1_N(_09909_),
    .A2_N(_09914_),
    .B1(_09909_),
    .B2(_09914_),
    .X(_09915_));
 sky130_fd_sc_hd__a2bb2o_2 _24259_ (.A1_N(_09908_),
    .A2_N(_09915_),
    .B1(_09908_),
    .B2(_09915_),
    .X(_09916_));
 sky130_fd_sc_hd__o2bb2ai_2 _24260_ (.A1_N(_09907_),
    .A2_N(_09916_),
    .B1(_09907_),
    .B2(_09916_),
    .Y(_09917_));
 sky130_fd_sc_hd__o22a_2 _24261_ (.A1(_09827_),
    .A2(_09828_),
    .B1(_09829_),
    .B2(_09839_),
    .X(_09918_));
 sky130_fd_sc_hd__o2bb2ai_2 _24262_ (.A1_N(_09917_),
    .A2_N(_09918_),
    .B1(_09917_),
    .B2(_09918_),
    .Y(_09919_));
 sky130_fd_sc_hd__buf_1 _24263_ (.A(_09766_),
    .X(_09920_));
 sky130_fd_sc_hd__o22a_2 _24264_ (.A1(_09846_),
    .A2(_09851_),
    .B1(_09920_),
    .B2(_09852_),
    .X(_09921_));
 sky130_fd_sc_hd__o22a_2 _24265_ (.A1(_09831_),
    .A2(_09837_),
    .B1(_09830_),
    .B2(_09838_),
    .X(_09922_));
 sky130_fd_sc_hd__o22a_2 _24266_ (.A1(_10588_),
    .A2(_09306_),
    .B1(_10588_),
    .B2(_09305_),
    .X(_09923_));
 sky130_fd_sc_hd__or4_2 _24267_ (.A(_10587_),
    .B(_09306_),
    .C(_10587_),
    .D(_09305_),
    .X(_09924_));
 sky130_fd_sc_hd__or2b_2 _24268_ (.A(_09923_),
    .B_N(_09924_),
    .X(_09925_));
 sky130_fd_sc_hd__o22a_2 _24269_ (.A1(_09773_),
    .A2(_09848_),
    .B1(_09310_),
    .B2(_09847_),
    .X(_09926_));
 sky130_fd_sc_hd__a2bb2oi_2 _24270_ (.A1_N(_09925_),
    .A2_N(_09926_),
    .B1(_09925_),
    .B2(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__a2bb2o_2 _24271_ (.A1_N(_09766_),
    .A2_N(_09927_),
    .B1(_09766_),
    .B2(_09927_),
    .X(_09928_));
 sky130_fd_sc_hd__a2bb2o_2 _24272_ (.A1_N(_09922_),
    .A2_N(_09928_),
    .B1(_09922_),
    .B2(_09928_),
    .X(_09929_));
 sky130_fd_sc_hd__a2bb2o_2 _24273_ (.A1_N(_09921_),
    .A2_N(_09929_),
    .B1(_09921_),
    .B2(_09929_),
    .X(_09930_));
 sky130_fd_sc_hd__o2bb2ai_2 _24274_ (.A1_N(_09919_),
    .A2_N(_09930_),
    .B1(_09919_),
    .B2(_09930_),
    .Y(_09931_));
 sky130_fd_sc_hd__o22a_2 _24275_ (.A1(_09840_),
    .A2(_09841_),
    .B1(_09842_),
    .B2(_09855_),
    .X(_09932_));
 sky130_fd_sc_hd__o2bb2a_2 _24276_ (.A1_N(_09931_),
    .A2_N(_09932_),
    .B1(_09931_),
    .B2(_09932_),
    .X(_09933_));
 sky130_vsdinv _24277_ (.A(_09933_),
    .Y(_09934_));
 sky130_fd_sc_hd__o21a_2 _24278_ (.A1(_09272_),
    .A2(_09865_),
    .B1(_09860_),
    .X(_09935_));
 sky130_fd_sc_hd__o22a_2 _24279_ (.A1(_09844_),
    .A2(_09853_),
    .B1(_09843_),
    .B2(_09854_),
    .X(_09936_));
 sky130_fd_sc_hd__a2bb2o_2 _24280_ (.A1_N(_09866_),
    .A2_N(_09936_),
    .B1(_09866_),
    .B2(_09936_),
    .X(_09937_));
 sky130_fd_sc_hd__a2bb2o_2 _24281_ (.A1_N(_09935_),
    .A2_N(_09937_),
    .B1(_09935_),
    .B2(_09937_),
    .X(_09938_));
 sky130_vsdinv _24282_ (.A(_09938_),
    .Y(_09939_));
 sky130_fd_sc_hd__a22o_2 _24283_ (.A1(_09934_),
    .A2(_09938_),
    .B1(_09933_),
    .B2(_09939_),
    .X(_09940_));
 sky130_fd_sc_hd__o22a_2 _24284_ (.A1(_09856_),
    .A2(_09857_),
    .B1(_09859_),
    .B2(_09868_),
    .X(_09941_));
 sky130_fd_sc_hd__a2bb2o_2 _24285_ (.A1_N(_09940_),
    .A2_N(_09941_),
    .B1(_09940_),
    .B2(_09941_),
    .X(_09942_));
 sky130_fd_sc_hd__o22a_2 _24286_ (.A1(_09862_),
    .A2(_09866_),
    .B1(_09861_),
    .B2(_09867_),
    .X(_09943_));
 sky130_fd_sc_hd__a2bb2o_2 _24287_ (.A1_N(_09472_),
    .A2_N(_09943_),
    .B1(_09472_),
    .B2(_09943_),
    .X(_09944_));
 sky130_fd_sc_hd__a2bb2o_2 _24288_ (.A1_N(_09630_),
    .A2_N(_09944_),
    .B1(_09630_),
    .B2(_09944_),
    .X(_09945_));
 sky130_fd_sc_hd__a2bb2o_2 _24289_ (.A1_N(_09942_),
    .A2_N(_09945_),
    .B1(_09942_),
    .B2(_09945_),
    .X(_09946_));
 sky130_fd_sc_hd__o22a_2 _24290_ (.A1(_09870_),
    .A2(_09871_),
    .B1(_09872_),
    .B2(_09875_),
    .X(_09947_));
 sky130_fd_sc_hd__a2bb2o_2 _24291_ (.A1_N(_09946_),
    .A2_N(_09947_),
    .B1(_09946_),
    .B2(_09947_),
    .X(_09948_));
 sky130_fd_sc_hd__o22a_2 _24292_ (.A1(_09563_),
    .A2(_09873_),
    .B1(_09564_),
    .B2(_09874_),
    .X(_09949_));
 sky130_fd_sc_hd__or2_2 _24293_ (.A(_09257_),
    .B(_09949_),
    .X(_09950_));
 sky130_fd_sc_hd__a21bo_2 _24294_ (.A1(_09719_),
    .A2(_09949_),
    .B1_N(_09950_),
    .X(_09951_));
 sky130_fd_sc_hd__a2bb2o_2 _24295_ (.A1_N(_09948_),
    .A2_N(_09951_),
    .B1(_09948_),
    .B2(_09951_),
    .X(_09952_));
 sky130_fd_sc_hd__o22a_2 _24296_ (.A1(_09876_),
    .A2(_09877_),
    .B1(_09878_),
    .B2(_09881_),
    .X(_09953_));
 sky130_fd_sc_hd__a2bb2o_2 _24297_ (.A1_N(_09952_),
    .A2_N(_09953_),
    .B1(_09952_),
    .B2(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__a2bb2o_2 _24298_ (.A1_N(_09880_),
    .A2_N(_09954_),
    .B1(_09880_),
    .B2(_09954_),
    .X(_09955_));
 sky130_fd_sc_hd__o22a_2 _24299_ (.A1(_09882_),
    .A2(_09883_),
    .B1(_09805_),
    .B2(_09884_),
    .X(_09956_));
 sky130_fd_sc_hd__and2_2 _24300_ (.A(_09955_),
    .B(_09956_),
    .X(_09957_));
 sky130_fd_sc_hd__or2_2 _24301_ (.A(_09955_),
    .B(_09956_),
    .X(_09958_));
 sky130_fd_sc_hd__or2b_2 _24302_ (.A(_09957_),
    .B_N(_09958_),
    .X(_09959_));
 sky130_fd_sc_hd__o21ai_2 _24303_ (.A1(_09888_),
    .A2(_09890_),
    .B1(_09887_),
    .Y(_09960_));
 sky130_fd_sc_hd__a2bb2o_2 _24304_ (.A1_N(_09959_),
    .A2_N(_09960_),
    .B1(_09959_),
    .B2(_09960_),
    .X(_02674_));
 sky130_fd_sc_hd__and4_2 _24305_ (.A(_09646_),
    .B(_06620_),
    .C(_11562_),
    .D(_11894_),
    .X(_09961_));
 sky130_fd_sc_hd__o22a_2 _24306_ (.A1(_10598_),
    .A2(_11896_),
    .B1(_09738_),
    .B2(_09429_),
    .X(_09962_));
 sky130_fd_sc_hd__nor2_2 _24307_ (.A(_09961_),
    .B(_09962_),
    .Y(_09963_));
 sky130_fd_sc_hd__nor2_2 _24308_ (.A(_09650_),
    .B(_09748_),
    .Y(_09964_));
 sky130_fd_sc_hd__a2bb2o_2 _24309_ (.A1_N(_09963_),
    .A2_N(_09964_),
    .B1(_09963_),
    .B2(_09964_),
    .X(_09965_));
 sky130_fd_sc_hd__a21oi_2 _24310_ (.A1(_09893_),
    .A2(_09894_),
    .B1(_09891_),
    .Y(_09966_));
 sky130_fd_sc_hd__o2bb2ai_2 _24311_ (.A1_N(_09965_),
    .A2_N(_09966_),
    .B1(_09965_),
    .B2(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__buf_1 _24312_ (.A(_09655_),
    .X(_09968_));
 sky130_fd_sc_hd__o22a_2 _24313_ (.A1(_09968_),
    .A2(_09311_),
    .B1(_09898_),
    .B2(_09902_),
    .X(_09969_));
 sky130_fd_sc_hd__and4_2 _24314_ (.A(_11569_),
    .B(_11886_),
    .C(_11573_),
    .D(_11883_),
    .X(_09970_));
 sky130_fd_sc_hd__nor2_2 _24315_ (.A(_09969_),
    .B(_09970_),
    .Y(_09971_));
 sky130_fd_sc_hd__buf_1 _24316_ (.A(_07289_),
    .X(_09972_));
 sky130_fd_sc_hd__nor2_2 _24317_ (.A(_09824_),
    .B(_09972_),
    .Y(_09973_));
 sky130_fd_sc_hd__a2bb2o_2 _24318_ (.A1_N(_09971_),
    .A2_N(_09973_),
    .B1(_09971_),
    .B2(_09973_),
    .X(_09974_));
 sky130_fd_sc_hd__o2bb2ai_2 _24319_ (.A1_N(_09967_),
    .A2_N(_09974_),
    .B1(_09967_),
    .B2(_09974_),
    .Y(_09975_));
 sky130_fd_sc_hd__o22a_2 _24320_ (.A1(_09895_),
    .A2(_09896_),
    .B1(_09897_),
    .B2(_09904_),
    .X(_09976_));
 sky130_fd_sc_hd__o2bb2ai_2 _24321_ (.A1_N(_09975_),
    .A2_N(_09976_),
    .B1(_09975_),
    .B2(_09976_),
    .Y(_09977_));
 sky130_fd_sc_hd__a21oi_2 _24322_ (.A1(_09912_),
    .A2(_09913_),
    .B1(_09911_),
    .Y(_09978_));
 sky130_fd_sc_hd__a21oi_2 _24323_ (.A1(_09901_),
    .A2(_09903_),
    .B1(_09900_),
    .Y(_09979_));
 sky130_fd_sc_hd__buf_1 _24324_ (.A(_09284_),
    .X(_09980_));
 sky130_fd_sc_hd__o22a_2 _24325_ (.A1(_09832_),
    .A2(_09302_),
    .B1(_06443_),
    .B2(_09699_),
    .X(_09981_));
 sky130_fd_sc_hd__and4_2 _24326_ (.A(_11577_),
    .B(_11879_),
    .C(_11582_),
    .D(_11875_),
    .X(_09982_));
 sky130_fd_sc_hd__or2_2 _24327_ (.A(_09981_),
    .B(_09982_),
    .X(_09983_));
 sky130_vsdinv _24328_ (.A(_09983_),
    .Y(_09984_));
 sky130_fd_sc_hd__or2_2 _24329_ (.A(_10588_),
    .B(_06275_),
    .X(_09985_));
 sky130_fd_sc_hd__a32o_2 _24330_ (.A1(_09980_),
    .A2(\pcpi_mul.rs2[24] ),
    .A3(_09984_),
    .B1(_09983_),
    .B2(_09985_),
    .X(_09986_));
 sky130_fd_sc_hd__a2bb2o_2 _24331_ (.A1_N(_09979_),
    .A2_N(_09986_),
    .B1(_09979_),
    .B2(_09986_),
    .X(_09987_));
 sky130_fd_sc_hd__a2bb2o_2 _24332_ (.A1_N(_09978_),
    .A2_N(_09987_),
    .B1(_09978_),
    .B2(_09987_),
    .X(_09988_));
 sky130_fd_sc_hd__o2bb2ai_2 _24333_ (.A1_N(_09977_),
    .A2_N(_09988_),
    .B1(_09977_),
    .B2(_09988_),
    .Y(_09989_));
 sky130_fd_sc_hd__o22a_2 _24334_ (.A1(_09905_),
    .A2(_09906_),
    .B1(_09907_),
    .B2(_09916_),
    .X(_09990_));
 sky130_fd_sc_hd__o2bb2ai_2 _24335_ (.A1_N(_09989_),
    .A2_N(_09990_),
    .B1(_09989_),
    .B2(_09990_),
    .Y(_09991_));
 sky130_fd_sc_hd__or2_2 _24336_ (.A(_09310_),
    .B(_09924_),
    .X(_09992_));
 sky130_fd_sc_hd__o21a_2 _24337_ (.A1(_09920_),
    .A2(_09927_),
    .B1(_09992_),
    .X(_09993_));
 sky130_fd_sc_hd__o22a_2 _24338_ (.A1(_09909_),
    .A2(_09914_),
    .B1(_09908_),
    .B2(_09915_),
    .X(_09994_));
 sky130_vsdinv _24339_ (.A(_09992_),
    .Y(_09995_));
 sky130_fd_sc_hd__and2_2 _24340_ (.A(_09772_),
    .B(_09923_),
    .X(_09996_));
 sky130_fd_sc_hd__or2_2 _24341_ (.A(_09995_),
    .B(_09996_),
    .X(_09997_));
 sky130_fd_sc_hd__a2bb2o_2 _24342_ (.A1_N(_09920_),
    .A2_N(_09997_),
    .B1(_09920_),
    .B2(_09997_),
    .X(_09998_));
 sky130_fd_sc_hd__a2bb2o_2 _24343_ (.A1_N(_09994_),
    .A2_N(_09998_),
    .B1(_09994_),
    .B2(_09998_),
    .X(_09999_));
 sky130_fd_sc_hd__a2bb2o_2 _24344_ (.A1_N(_09993_),
    .A2_N(_09999_),
    .B1(_09993_),
    .B2(_09999_),
    .X(_10000_));
 sky130_fd_sc_hd__o2bb2ai_2 _24345_ (.A1_N(_09991_),
    .A2_N(_10000_),
    .B1(_09991_),
    .B2(_10000_),
    .Y(_10001_));
 sky130_fd_sc_hd__o22a_2 _24346_ (.A1(_09917_),
    .A2(_09918_),
    .B1(_09919_),
    .B2(_09930_),
    .X(_10002_));
 sky130_fd_sc_hd__o2bb2a_2 _24347_ (.A1_N(_10001_),
    .A2_N(_10002_),
    .B1(_10001_),
    .B2(_10002_),
    .X(_10003_));
 sky130_vsdinv _24348_ (.A(_10003_),
    .Y(_10004_));
 sky130_fd_sc_hd__buf_1 _24349_ (.A(_09935_),
    .X(_10005_));
 sky130_fd_sc_hd__buf_1 _24350_ (.A(_10005_),
    .X(_10006_));
 sky130_fd_sc_hd__buf_1 _24351_ (.A(_09866_),
    .X(_10007_));
 sky130_fd_sc_hd__buf_1 _24352_ (.A(_10007_),
    .X(_10008_));
 sky130_fd_sc_hd__o22a_2 _24353_ (.A1(_09922_),
    .A2(_09928_),
    .B1(_09921_),
    .B2(_09929_),
    .X(_10009_));
 sky130_fd_sc_hd__a2bb2o_2 _24354_ (.A1_N(_10008_),
    .A2_N(_10009_),
    .B1(_10007_),
    .B2(_10009_),
    .X(_10010_));
 sky130_fd_sc_hd__a2bb2o_2 _24355_ (.A1_N(_10006_),
    .A2_N(_10010_),
    .B1(_10006_),
    .B2(_10010_),
    .X(_10011_));
 sky130_vsdinv _24356_ (.A(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__a22o_2 _24357_ (.A1(_10004_),
    .A2(_10011_),
    .B1(_10003_),
    .B2(_10012_),
    .X(_10013_));
 sky130_fd_sc_hd__o22a_2 _24358_ (.A1(_09931_),
    .A2(_09932_),
    .B1(_09934_),
    .B2(_09938_),
    .X(_10014_));
 sky130_fd_sc_hd__a2bb2o_2 _24359_ (.A1_N(_10013_),
    .A2_N(_10014_),
    .B1(_10013_),
    .B2(_10014_),
    .X(_10015_));
 sky130_fd_sc_hd__buf_1 _24360_ (.A(_09630_),
    .X(_10016_));
 sky130_fd_sc_hd__buf_1 _24361_ (.A(_09563_),
    .X(_10017_));
 sky130_fd_sc_hd__buf_1 _24362_ (.A(_10008_),
    .X(_10018_));
 sky130_fd_sc_hd__o22a_2 _24363_ (.A1(_10018_),
    .A2(_09936_),
    .B1(_10006_),
    .B2(_09937_),
    .X(_10019_));
 sky130_fd_sc_hd__a2bb2o_2 _24364_ (.A1_N(_10017_),
    .A2_N(_10019_),
    .B1(_10017_),
    .B2(_10019_),
    .X(_10020_));
 sky130_fd_sc_hd__a2bb2o_2 _24365_ (.A1_N(_10016_),
    .A2_N(_10020_),
    .B1(_10016_),
    .B2(_10020_),
    .X(_10021_));
 sky130_fd_sc_hd__a2bb2o_2 _24366_ (.A1_N(_10015_),
    .A2_N(_10021_),
    .B1(_10015_),
    .B2(_10021_),
    .X(_10022_));
 sky130_fd_sc_hd__o22a_2 _24367_ (.A1(_09940_),
    .A2(_09941_),
    .B1(_09942_),
    .B2(_09945_),
    .X(_10023_));
 sky130_fd_sc_hd__a2bb2o_2 _24368_ (.A1_N(_10022_),
    .A2_N(_10023_),
    .B1(_10022_),
    .B2(_10023_),
    .X(_10024_));
 sky130_fd_sc_hd__buf_1 _24369_ (.A(_09719_),
    .X(_10025_));
 sky130_fd_sc_hd__buf_1 _24370_ (.A(_09563_),
    .X(_10026_));
 sky130_fd_sc_hd__buf_1 _24371_ (.A(_10026_),
    .X(_10027_));
 sky130_fd_sc_hd__buf_1 _24372_ (.A(_09630_),
    .X(_10028_));
 sky130_fd_sc_hd__o22a_2 _24373_ (.A1(_10027_),
    .A2(_09943_),
    .B1(_10028_),
    .B2(_09944_),
    .X(_10029_));
 sky130_fd_sc_hd__or2_2 _24374_ (.A(_10025_),
    .B(_10029_),
    .X(_10030_));
 sky130_fd_sc_hd__a21bo_2 _24375_ (.A1(_10025_),
    .A2(_10029_),
    .B1_N(_10030_),
    .X(_10031_));
 sky130_fd_sc_hd__a2bb2o_2 _24376_ (.A1_N(_10024_),
    .A2_N(_10031_),
    .B1(_10024_),
    .B2(_10031_),
    .X(_10032_));
 sky130_fd_sc_hd__o22a_2 _24377_ (.A1(_09946_),
    .A2(_09947_),
    .B1(_09948_),
    .B2(_09951_),
    .X(_10033_));
 sky130_fd_sc_hd__a2bb2o_2 _24378_ (.A1_N(_10032_),
    .A2_N(_10033_),
    .B1(_10032_),
    .B2(_10033_),
    .X(_10034_));
 sky130_fd_sc_hd__a2bb2o_2 _24379_ (.A1_N(_09950_),
    .A2_N(_10034_),
    .B1(_09950_),
    .B2(_10034_),
    .X(_10035_));
 sky130_fd_sc_hd__o22a_2 _24380_ (.A1(_09952_),
    .A2(_09953_),
    .B1(_09880_),
    .B2(_09954_),
    .X(_10036_));
 sky130_fd_sc_hd__or2_2 _24381_ (.A(_10035_),
    .B(_10036_),
    .X(_10037_));
 sky130_fd_sc_hd__a21bo_2 _24382_ (.A1(_10035_),
    .A2(_10036_),
    .B1_N(_10037_),
    .X(_10038_));
 sky130_fd_sc_hd__or2_2 _24383_ (.A(_09888_),
    .B(_09959_),
    .X(_10039_));
 sky130_fd_sc_hd__or3_2 _24384_ (.A(_09729_),
    .B(_09813_),
    .C(_10039_),
    .X(_10040_));
 sky130_fd_sc_hd__or2_2 _24385_ (.A(_09731_),
    .B(_10040_),
    .X(_10041_));
 sky130_fd_sc_hd__o221a_2 _24386_ (.A1(_09887_),
    .A2(_09957_),
    .B1(_09889_),
    .B2(_10039_),
    .C1(_09958_),
    .X(_10042_));
 sky130_fd_sc_hd__o221a_2 _24387_ (.A1(_09732_),
    .A2(_10040_),
    .B1(_09372_),
    .B2(_10041_),
    .C1(_10042_),
    .X(_10043_));
 sky130_fd_sc_hd__a2bb2oi_2 _24388_ (.A1_N(_10038_),
    .A2_N(_10043_),
    .B1(_10038_),
    .B2(_10043_),
    .Y(_02675_));
 sky130_fd_sc_hd__buf_1 _24389_ (.A(_09646_),
    .X(_10044_));
 sky130_fd_sc_hd__and4_2 _24390_ (.A(_10044_),
    .B(_09429_),
    .C(_11563_),
    .D(_11890_),
    .X(_10045_));
 sky130_fd_sc_hd__buf_1 _24391_ (.A(_09738_),
    .X(_10046_));
 sky130_fd_sc_hd__o22a_2 _24392_ (.A1(_10599_),
    .A2(_11894_),
    .B1(_10046_),
    .B2(_09748_),
    .X(_10047_));
 sky130_fd_sc_hd__nor2_2 _24393_ (.A(_10045_),
    .B(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__buf_1 _24394_ (.A(_09650_),
    .X(_10049_));
 sky130_fd_sc_hd__nor2_2 _24395_ (.A(_10049_),
    .B(_09311_),
    .Y(_10050_));
 sky130_fd_sc_hd__a2bb2o_2 _24396_ (.A1_N(_10048_),
    .A2_N(_10050_),
    .B1(_10048_),
    .B2(_10050_),
    .X(_10051_));
 sky130_fd_sc_hd__a21oi_2 _24397_ (.A1(_09963_),
    .A2(_09964_),
    .B1(_09961_),
    .Y(_10052_));
 sky130_fd_sc_hd__o2bb2ai_2 _24398_ (.A1_N(_10051_),
    .A2_N(_10052_),
    .B1(_10051_),
    .B2(_10052_),
    .Y(_10053_));
 sky130_fd_sc_hd__o22a_2 _24399_ (.A1(_09968_),
    .A2(_09902_),
    .B1(_09898_),
    .B2(_09972_),
    .X(_10054_));
 sky130_fd_sc_hd__and4_2 _24400_ (.A(_11569_),
    .B(_11883_),
    .C(_11573_),
    .D(_11881_),
    .X(_10055_));
 sky130_fd_sc_hd__nor2_2 _24401_ (.A(_10054_),
    .B(_10055_),
    .Y(_10056_));
 sky130_fd_sc_hd__buf_1 _24402_ (.A(_09302_),
    .X(_10057_));
 sky130_fd_sc_hd__nor2_2 _24403_ (.A(_09824_),
    .B(_10057_),
    .Y(_10058_));
 sky130_fd_sc_hd__a2bb2o_2 _24404_ (.A1_N(_10056_),
    .A2_N(_10058_),
    .B1(_10056_),
    .B2(_10058_),
    .X(_10059_));
 sky130_fd_sc_hd__o2bb2ai_2 _24405_ (.A1_N(_10053_),
    .A2_N(_10059_),
    .B1(_10053_),
    .B2(_10059_),
    .Y(_10060_));
 sky130_fd_sc_hd__o22a_2 _24406_ (.A1(_09965_),
    .A2(_09966_),
    .B1(_09967_),
    .B2(_09974_),
    .X(_10061_));
 sky130_fd_sc_hd__o2bb2ai_2 _24407_ (.A1_N(_10060_),
    .A2_N(_10061_),
    .B1(_10060_),
    .B2(_10061_),
    .Y(_10062_));
 sky130_fd_sc_hd__buf_1 _24408_ (.A(_09985_),
    .X(_10063_));
 sky130_fd_sc_hd__o21ba_2 _24409_ (.A1(_09983_),
    .A2(_10063_),
    .B1_N(_09982_),
    .X(_10064_));
 sky130_fd_sc_hd__a21oi_2 _24410_ (.A1(_09971_),
    .A2(_09973_),
    .B1(_09970_),
    .Y(_10065_));
 sky130_fd_sc_hd__buf_1 _24411_ (.A(_09699_),
    .X(_10066_));
 sky130_fd_sc_hd__nor2_2 _24412_ (.A(_09832_),
    .B(_10066_),
    .Y(_10067_));
 sky130_fd_sc_hd__or2_2 _24413_ (.A(_10588_),
    .B(_06443_),
    .X(_10068_));
 sky130_vsdinv _24414_ (.A(_10068_),
    .Y(_10069_));
 sky130_fd_sc_hd__a2bb2o_2 _24415_ (.A1_N(_10067_),
    .A2_N(_10069_),
    .B1(_10067_),
    .B2(_10069_),
    .X(_10070_));
 sky130_fd_sc_hd__a2bb2o_2 _24416_ (.A1_N(_10063_),
    .A2_N(_10070_),
    .B1(_09985_),
    .B2(_10070_),
    .X(_10071_));
 sky130_fd_sc_hd__a2bb2o_2 _24417_ (.A1_N(_10065_),
    .A2_N(_10071_),
    .B1(_10065_),
    .B2(_10071_),
    .X(_10072_));
 sky130_fd_sc_hd__a2bb2o_2 _24418_ (.A1_N(_10064_),
    .A2_N(_10072_),
    .B1(_10064_),
    .B2(_10072_),
    .X(_10073_));
 sky130_fd_sc_hd__o2bb2ai_2 _24419_ (.A1_N(_10062_),
    .A2_N(_10073_),
    .B1(_10062_),
    .B2(_10073_),
    .Y(_10074_));
 sky130_fd_sc_hd__o22a_2 _24420_ (.A1(_09975_),
    .A2(_09976_),
    .B1(_09977_),
    .B2(_09988_),
    .X(_10075_));
 sky130_fd_sc_hd__o2bb2ai_2 _24421_ (.A1_N(_10074_),
    .A2_N(_10075_),
    .B1(_10074_),
    .B2(_10075_),
    .Y(_10076_));
 sky130_fd_sc_hd__o21a_2 _24422_ (.A1(_09920_),
    .A2(_09997_),
    .B1(_09992_),
    .X(_10077_));
 sky130_fd_sc_hd__buf_1 _24423_ (.A(_10077_),
    .X(_10078_));
 sky130_fd_sc_hd__o22a_2 _24424_ (.A1(_09979_),
    .A2(_09986_),
    .B1(_09978_),
    .B2(_09987_),
    .X(_10079_));
 sky130_fd_sc_hd__a2bb2o_2 _24425_ (.A1_N(_09998_),
    .A2_N(_10079_),
    .B1(_09998_),
    .B2(_10079_),
    .X(_10080_));
 sky130_fd_sc_hd__a2bb2o_2 _24426_ (.A1_N(_10078_),
    .A2_N(_10080_),
    .B1(_10078_),
    .B2(_10080_),
    .X(_10081_));
 sky130_fd_sc_hd__o2bb2ai_2 _24427_ (.A1_N(_10076_),
    .A2_N(_10081_),
    .B1(_10076_),
    .B2(_10081_),
    .Y(_10082_));
 sky130_fd_sc_hd__o22a_2 _24428_ (.A1(_09989_),
    .A2(_09990_),
    .B1(_09991_),
    .B2(_10000_),
    .X(_10083_));
 sky130_fd_sc_hd__o2bb2a_2 _24429_ (.A1_N(_10082_),
    .A2_N(_10083_),
    .B1(_10082_),
    .B2(_10083_),
    .X(_10084_));
 sky130_vsdinv _24430_ (.A(_10084_),
    .Y(_10085_));
 sky130_fd_sc_hd__buf_1 _24431_ (.A(_09998_),
    .X(_10086_));
 sky130_fd_sc_hd__buf_1 _24432_ (.A(_10086_),
    .X(_10087_));
 sky130_fd_sc_hd__o22a_2 _24433_ (.A1(_09994_),
    .A2(_10087_),
    .B1(_09993_),
    .B2(_09999_),
    .X(_10088_));
 sky130_fd_sc_hd__a2bb2o_2 _24434_ (.A1_N(_10007_),
    .A2_N(_10088_),
    .B1(_10007_),
    .B2(_10088_),
    .X(_10089_));
 sky130_fd_sc_hd__a2bb2o_2 _24435_ (.A1_N(_10005_),
    .A2_N(_10089_),
    .B1(_10005_),
    .B2(_10089_),
    .X(_10090_));
 sky130_vsdinv _24436_ (.A(_10090_),
    .Y(_10091_));
 sky130_fd_sc_hd__a22o_2 _24437_ (.A1(_10085_),
    .A2(_10090_),
    .B1(_10084_),
    .B2(_10091_),
    .X(_10092_));
 sky130_fd_sc_hd__o22a_2 _24438_ (.A1(_10001_),
    .A2(_10002_),
    .B1(_10004_),
    .B2(_10011_),
    .X(_10093_));
 sky130_fd_sc_hd__a2bb2o_2 _24439_ (.A1_N(_10092_),
    .A2_N(_10093_),
    .B1(_10092_),
    .B2(_10093_),
    .X(_10094_));
 sky130_fd_sc_hd__o22a_2 _24440_ (.A1(_10008_),
    .A2(_10009_),
    .B1(_10006_),
    .B2(_10010_),
    .X(_10095_));
 sky130_fd_sc_hd__a2bb2o_2 _24441_ (.A1_N(_10017_),
    .A2_N(_10095_),
    .B1(_10017_),
    .B2(_10095_),
    .X(_10096_));
 sky130_fd_sc_hd__a2bb2o_2 _24442_ (.A1_N(_10016_),
    .A2_N(_10096_),
    .B1(_10016_),
    .B2(_10096_),
    .X(_10097_));
 sky130_fd_sc_hd__a2bb2o_2 _24443_ (.A1_N(_10094_),
    .A2_N(_10097_),
    .B1(_10094_),
    .B2(_10097_),
    .X(_10098_));
 sky130_fd_sc_hd__o22a_2 _24444_ (.A1(_10013_),
    .A2(_10014_),
    .B1(_10015_),
    .B2(_10021_),
    .X(_10099_));
 sky130_fd_sc_hd__a2bb2o_2 _24445_ (.A1_N(_10098_),
    .A2_N(_10099_),
    .B1(_10098_),
    .B2(_10099_),
    .X(_10100_));
 sky130_fd_sc_hd__o22a_2 _24446_ (.A1(_10026_),
    .A2(_10019_),
    .B1(_10028_),
    .B2(_10020_),
    .X(_10101_));
 sky130_fd_sc_hd__or2_2 _24447_ (.A(_09719_),
    .B(_10101_),
    .X(_10102_));
 sky130_fd_sc_hd__a21bo_2 _24448_ (.A1(_10025_),
    .A2(_10101_),
    .B1_N(_10102_),
    .X(_10103_));
 sky130_fd_sc_hd__a2bb2o_2 _24449_ (.A1_N(_10100_),
    .A2_N(_10103_),
    .B1(_10100_),
    .B2(_10103_),
    .X(_10104_));
 sky130_fd_sc_hd__o22a_2 _24450_ (.A1(_10022_),
    .A2(_10023_),
    .B1(_10024_),
    .B2(_10031_),
    .X(_10105_));
 sky130_fd_sc_hd__a2bb2o_2 _24451_ (.A1_N(_10104_),
    .A2_N(_10105_),
    .B1(_10104_),
    .B2(_10105_),
    .X(_10106_));
 sky130_fd_sc_hd__a2bb2o_2 _24452_ (.A1_N(_10030_),
    .A2_N(_10106_),
    .B1(_10030_),
    .B2(_10106_),
    .X(_10107_));
 sky130_fd_sc_hd__o22a_2 _24453_ (.A1(_10032_),
    .A2(_10033_),
    .B1(_09950_),
    .B2(_10034_),
    .X(_10108_));
 sky130_fd_sc_hd__or2_2 _24454_ (.A(_10107_),
    .B(_10108_),
    .X(_10109_));
 sky130_fd_sc_hd__a21bo_2 _24455_ (.A1(_10107_),
    .A2(_10108_),
    .B1_N(_10109_),
    .X(_10110_));
 sky130_fd_sc_hd__o21ai_2 _24456_ (.A1(_10038_),
    .A2(_10043_),
    .B1(_10037_),
    .Y(_10111_));
 sky130_fd_sc_hd__a2bb2o_2 _24457_ (.A1_N(_10110_),
    .A2_N(_10111_),
    .B1(_10110_),
    .B2(_10111_),
    .X(_02676_));
 sky130_fd_sc_hd__and4_2 _24458_ (.A(_10044_),
    .B(_09748_),
    .C(_11563_),
    .D(_11886_),
    .X(_10112_));
 sky130_fd_sc_hd__o22a_2 _24459_ (.A1(_10599_),
    .A2(_11890_),
    .B1(_10046_),
    .B2(_09311_),
    .X(_10113_));
 sky130_fd_sc_hd__nor2_2 _24460_ (.A(_10112_),
    .B(_10113_),
    .Y(_10114_));
 sky130_fd_sc_hd__nor2_2 _24461_ (.A(_10049_),
    .B(_09902_),
    .Y(_10115_));
 sky130_fd_sc_hd__a2bb2o_2 _24462_ (.A1_N(_10114_),
    .A2_N(_10115_),
    .B1(_10114_),
    .B2(_10115_),
    .X(_10116_));
 sky130_fd_sc_hd__a21oi_2 _24463_ (.A1(_10048_),
    .A2(_10050_),
    .B1(_10045_),
    .Y(_10117_));
 sky130_fd_sc_hd__o2bb2ai_2 _24464_ (.A1_N(_10116_),
    .A2_N(_10117_),
    .B1(_10116_),
    .B2(_10117_),
    .Y(_10118_));
 sky130_fd_sc_hd__o22a_2 _24465_ (.A1(_09968_),
    .A2(_09972_),
    .B1(_09898_),
    .B2(_10057_),
    .X(_10119_));
 sky130_fd_sc_hd__and4_2 _24466_ (.A(_11569_),
    .B(_11881_),
    .C(_11573_),
    .D(_11879_),
    .X(_10120_));
 sky130_fd_sc_hd__nor2_2 _24467_ (.A(_10119_),
    .B(_10120_),
    .Y(_10121_));
 sky130_fd_sc_hd__nor2_2 _24468_ (.A(_09824_),
    .B(_10066_),
    .Y(_10122_));
 sky130_fd_sc_hd__a2bb2o_2 _24469_ (.A1_N(_10121_),
    .A2_N(_10122_),
    .B1(_10121_),
    .B2(_10122_),
    .X(_10123_));
 sky130_fd_sc_hd__o2bb2ai_2 _24470_ (.A1_N(_10118_),
    .A2_N(_10123_),
    .B1(_10118_),
    .B2(_10123_),
    .Y(_10124_));
 sky130_fd_sc_hd__o22a_2 _24471_ (.A1(_10051_),
    .A2(_10052_),
    .B1(_10053_),
    .B2(_10059_),
    .X(_10125_));
 sky130_fd_sc_hd__o2bb2ai_2 _24472_ (.A1_N(_10124_),
    .A2_N(_10125_),
    .B1(_10124_),
    .B2(_10125_),
    .Y(_10126_));
 sky130_fd_sc_hd__o32a_2 _24473_ (.A1(_09832_),
    .A2(_10066_),
    .A3(_10068_),
    .B1(_10063_),
    .B2(_10070_),
    .X(_10127_));
 sky130_fd_sc_hd__a21oi_2 _24474_ (.A1(_10056_),
    .A2(_10058_),
    .B1(_10055_),
    .Y(_10128_));
 sky130_fd_sc_hd__or2_2 _24475_ (.A(_10588_),
    .B(_09832_),
    .X(_10129_));
 sky130_fd_sc_hd__a32o_2 _24476_ (.A1(_09284_),
    .A2(_11577_),
    .A3(_10069_),
    .B1(_10068_),
    .B2(_10129_),
    .X(_10130_));
 sky130_fd_sc_hd__a2bb2o_2 _24477_ (.A1_N(_10063_),
    .A2_N(_10130_),
    .B1(_10063_),
    .B2(_10130_),
    .X(_10131_));
 sky130_fd_sc_hd__a2bb2o_2 _24478_ (.A1_N(_10128_),
    .A2_N(_10131_),
    .B1(_10128_),
    .B2(_10131_),
    .X(_10132_));
 sky130_fd_sc_hd__a2bb2o_2 _24479_ (.A1_N(_10127_),
    .A2_N(_10132_),
    .B1(_10127_),
    .B2(_10132_),
    .X(_10133_));
 sky130_fd_sc_hd__o2bb2ai_2 _24480_ (.A1_N(_10126_),
    .A2_N(_10133_),
    .B1(_10126_),
    .B2(_10133_),
    .Y(_10134_));
 sky130_fd_sc_hd__o22a_2 _24481_ (.A1(_10060_),
    .A2(_10061_),
    .B1(_10062_),
    .B2(_10073_),
    .X(_10135_));
 sky130_fd_sc_hd__o2bb2ai_2 _24482_ (.A1_N(_10134_),
    .A2_N(_10135_),
    .B1(_10134_),
    .B2(_10135_),
    .Y(_10136_));
 sky130_fd_sc_hd__o22a_2 _24483_ (.A1(_10065_),
    .A2(_10071_),
    .B1(_10064_),
    .B2(_10072_),
    .X(_10137_));
 sky130_fd_sc_hd__a2bb2o_2 _24484_ (.A1_N(_10086_),
    .A2_N(_10137_),
    .B1(_10086_),
    .B2(_10137_),
    .X(_10138_));
 sky130_fd_sc_hd__a2bb2o_2 _24485_ (.A1_N(_10078_),
    .A2_N(_10138_),
    .B1(_10078_),
    .B2(_10138_),
    .X(_10139_));
 sky130_fd_sc_hd__o2bb2ai_2 _24486_ (.A1_N(_10136_),
    .A2_N(_10139_),
    .B1(_10136_),
    .B2(_10139_),
    .Y(_10140_));
 sky130_fd_sc_hd__o22a_2 _24487_ (.A1(_10074_),
    .A2(_10075_),
    .B1(_10076_),
    .B2(_10081_),
    .X(_10141_));
 sky130_fd_sc_hd__o2bb2a_2 _24488_ (.A1_N(_10140_),
    .A2_N(_10141_),
    .B1(_10140_),
    .B2(_10141_),
    .X(_10142_));
 sky130_vsdinv _24489_ (.A(_10142_),
    .Y(_10143_));
 sky130_fd_sc_hd__o22a_2 _24490_ (.A1(_10086_),
    .A2(_10079_),
    .B1(_10078_),
    .B2(_10080_),
    .X(_10144_));
 sky130_fd_sc_hd__a2bb2o_2 _24491_ (.A1_N(_10007_),
    .A2_N(_10144_),
    .B1(_10007_),
    .B2(_10144_),
    .X(_10145_));
 sky130_fd_sc_hd__a2bb2o_2 _24492_ (.A1_N(_10005_),
    .A2_N(_10145_),
    .B1(_10005_),
    .B2(_10145_),
    .X(_10146_));
 sky130_vsdinv _24493_ (.A(_10146_),
    .Y(_10147_));
 sky130_fd_sc_hd__a22o_2 _24494_ (.A1(_10143_),
    .A2(_10146_),
    .B1(_10142_),
    .B2(_10147_),
    .X(_10148_));
 sky130_fd_sc_hd__o22a_2 _24495_ (.A1(_10082_),
    .A2(_10083_),
    .B1(_10085_),
    .B2(_10090_),
    .X(_10149_));
 sky130_fd_sc_hd__a2bb2o_2 _24496_ (.A1_N(_10148_),
    .A2_N(_10149_),
    .B1(_10148_),
    .B2(_10149_),
    .X(_10150_));
 sky130_fd_sc_hd__buf_1 _24497_ (.A(_10005_),
    .X(_10151_));
 sky130_fd_sc_hd__o22a_2 _24498_ (.A1(_10018_),
    .A2(_10088_),
    .B1(_10151_),
    .B2(_10089_),
    .X(_10152_));
 sky130_fd_sc_hd__a2bb2o_2 _24499_ (.A1_N(_10017_),
    .A2_N(_10152_),
    .B1(_10017_),
    .B2(_10152_),
    .X(_10153_));
 sky130_fd_sc_hd__a2bb2o_2 _24500_ (.A1_N(_10016_),
    .A2_N(_10153_),
    .B1(_10028_),
    .B2(_10153_),
    .X(_10154_));
 sky130_fd_sc_hd__a2bb2o_2 _24501_ (.A1_N(_10150_),
    .A2_N(_10154_),
    .B1(_10150_),
    .B2(_10154_),
    .X(_10155_));
 sky130_fd_sc_hd__o22a_2 _24502_ (.A1(_10092_),
    .A2(_10093_),
    .B1(_10094_),
    .B2(_10097_),
    .X(_10156_));
 sky130_fd_sc_hd__a2bb2o_2 _24503_ (.A1_N(_10155_),
    .A2_N(_10156_),
    .B1(_10155_),
    .B2(_10156_),
    .X(_10157_));
 sky130_fd_sc_hd__o22a_2 _24504_ (.A1(_10026_),
    .A2(_10095_),
    .B1(_10028_),
    .B2(_10096_),
    .X(_10158_));
 sky130_fd_sc_hd__or2_2 _24505_ (.A(_09719_),
    .B(_10158_),
    .X(_10159_));
 sky130_fd_sc_hd__a21bo_2 _24506_ (.A1(_10025_),
    .A2(_10158_),
    .B1_N(_10159_),
    .X(_10160_));
 sky130_fd_sc_hd__a2bb2o_2 _24507_ (.A1_N(_10157_),
    .A2_N(_10160_),
    .B1(_10157_),
    .B2(_10160_),
    .X(_10161_));
 sky130_fd_sc_hd__o22a_2 _24508_ (.A1(_10098_),
    .A2(_10099_),
    .B1(_10100_),
    .B2(_10103_),
    .X(_10162_));
 sky130_fd_sc_hd__a2bb2o_2 _24509_ (.A1_N(_10161_),
    .A2_N(_10162_),
    .B1(_10161_),
    .B2(_10162_),
    .X(_10163_));
 sky130_fd_sc_hd__a2bb2o_2 _24510_ (.A1_N(_10102_),
    .A2_N(_10163_),
    .B1(_10102_),
    .B2(_10163_),
    .X(_10164_));
 sky130_fd_sc_hd__o22a_2 _24511_ (.A1(_10104_),
    .A2(_10105_),
    .B1(_10030_),
    .B2(_10106_),
    .X(_10165_));
 sky130_fd_sc_hd__or2_2 _24512_ (.A(_10164_),
    .B(_10165_),
    .X(_10166_));
 sky130_fd_sc_hd__a21bo_2 _24513_ (.A1(_10164_),
    .A2(_10165_),
    .B1_N(_10166_),
    .X(_10167_));
 sky130_fd_sc_hd__a22o_2 _24514_ (.A1(_10107_),
    .A2(_10108_),
    .B1(_10037_),
    .B2(_10109_),
    .X(_10168_));
 sky130_fd_sc_hd__o31a_2 _24515_ (.A1(_10038_),
    .A2(_10110_),
    .A3(_10043_),
    .B1(_10168_),
    .X(_10169_));
 sky130_fd_sc_hd__a2bb2oi_2 _24516_ (.A1_N(_10167_),
    .A2_N(_10169_),
    .B1(_10167_),
    .B2(_10169_),
    .Y(_02677_));
 sky130_fd_sc_hd__and4_2 _24517_ (.A(_10044_),
    .B(_09311_),
    .C(_11563_),
    .D(_11883_),
    .X(_10170_));
 sky130_fd_sc_hd__o22a_2 _24518_ (.A1(_10599_),
    .A2(_11886_),
    .B1(_10046_),
    .B2(_09902_),
    .X(_10171_));
 sky130_fd_sc_hd__nor2_2 _24519_ (.A(_10170_),
    .B(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__nor2_2 _24520_ (.A(_10049_),
    .B(_09972_),
    .Y(_10173_));
 sky130_fd_sc_hd__a2bb2o_2 _24521_ (.A1_N(_10172_),
    .A2_N(_10173_),
    .B1(_10172_),
    .B2(_10173_),
    .X(_10174_));
 sky130_fd_sc_hd__a21oi_2 _24522_ (.A1(_10114_),
    .A2(_10115_),
    .B1(_10112_),
    .Y(_10175_));
 sky130_fd_sc_hd__o2bb2ai_2 _24523_ (.A1_N(_10174_),
    .A2_N(_10175_),
    .B1(_10174_),
    .B2(_10175_),
    .Y(_10176_));
 sky130_fd_sc_hd__o22a_2 _24524_ (.A1(_09655_),
    .A2(_10057_),
    .B1(_09898_),
    .B2(_09699_),
    .X(_10177_));
 sky130_fd_sc_hd__and4_2 _24525_ (.A(_11569_),
    .B(_11879_),
    .C(_11573_),
    .D(_11875_),
    .X(_10178_));
 sky130_fd_sc_hd__or2_2 _24526_ (.A(_10177_),
    .B(_10178_),
    .X(_10179_));
 sky130_vsdinv _24527_ (.A(_10179_),
    .Y(_10180_));
 sky130_fd_sc_hd__or2_2 _24528_ (.A(_10589_),
    .B(_09824_),
    .X(_10181_));
 sky130_fd_sc_hd__a32o_2 _24529_ (.A1(_09980_),
    .A2(\pcpi_mul.rs2[27] ),
    .A3(_10180_),
    .B1(_10179_),
    .B2(_10181_),
    .X(_10182_));
 sky130_fd_sc_hd__o2bb2ai_2 _24530_ (.A1_N(_10176_),
    .A2_N(_10182_),
    .B1(_10176_),
    .B2(_10182_),
    .Y(_10183_));
 sky130_fd_sc_hd__o22a_2 _24531_ (.A1(_10116_),
    .A2(_10117_),
    .B1(_10118_),
    .B2(_10123_),
    .X(_10184_));
 sky130_fd_sc_hd__o2bb2ai_2 _24532_ (.A1_N(_10183_),
    .A2_N(_10184_),
    .B1(_10183_),
    .B2(_10184_),
    .Y(_10185_));
 sky130_fd_sc_hd__o22a_2 _24533_ (.A1(_10068_),
    .A2(_10129_),
    .B1(_10063_),
    .B2(_10130_),
    .X(_10186_));
 sky130_fd_sc_hd__buf_1 _24534_ (.A(_10186_),
    .X(_10187_));
 sky130_fd_sc_hd__a21oi_2 _24535_ (.A1(_10121_),
    .A2(_10122_),
    .B1(_10120_),
    .Y(_10188_));
 sky130_fd_sc_hd__a2bb2o_2 _24536_ (.A1_N(_10131_),
    .A2_N(_10188_),
    .B1(_10131_),
    .B2(_10188_),
    .X(_10189_));
 sky130_fd_sc_hd__a2bb2o_2 _24537_ (.A1_N(_10187_),
    .A2_N(_10189_),
    .B1(_10186_),
    .B2(_10189_),
    .X(_10190_));
 sky130_fd_sc_hd__o2bb2ai_2 _24538_ (.A1_N(_10185_),
    .A2_N(_10190_),
    .B1(_10185_),
    .B2(_10190_),
    .Y(_10191_));
 sky130_fd_sc_hd__o22a_2 _24539_ (.A1(_10124_),
    .A2(_10125_),
    .B1(_10126_),
    .B2(_10133_),
    .X(_10192_));
 sky130_fd_sc_hd__o2bb2ai_2 _24540_ (.A1_N(_10191_),
    .A2_N(_10192_),
    .B1(_10191_),
    .B2(_10192_),
    .Y(_10193_));
 sky130_fd_sc_hd__buf_1 _24541_ (.A(_10077_),
    .X(_10194_));
 sky130_fd_sc_hd__buf_1 _24542_ (.A(_10131_),
    .X(_10195_));
 sky130_fd_sc_hd__o22a_2 _24543_ (.A1(_10128_),
    .A2(_10195_),
    .B1(_10127_),
    .B2(_10132_),
    .X(_10196_));
 sky130_fd_sc_hd__a2bb2o_2 _24544_ (.A1_N(_10086_),
    .A2_N(_10196_),
    .B1(_10086_),
    .B2(_10196_),
    .X(_10197_));
 sky130_fd_sc_hd__a2bb2o_2 _24545_ (.A1_N(_10194_),
    .A2_N(_10197_),
    .B1(_10194_),
    .B2(_10197_),
    .X(_10198_));
 sky130_fd_sc_hd__o2bb2ai_2 _24546_ (.A1_N(_10193_),
    .A2_N(_10198_),
    .B1(_10193_),
    .B2(_10198_),
    .Y(_10199_));
 sky130_fd_sc_hd__o22a_2 _24547_ (.A1(_10134_),
    .A2(_10135_),
    .B1(_10136_),
    .B2(_10139_),
    .X(_10200_));
 sky130_fd_sc_hd__o2bb2a_2 _24548_ (.A1_N(_10199_),
    .A2_N(_10200_),
    .B1(_10199_),
    .B2(_10200_),
    .X(_10201_));
 sky130_vsdinv _24549_ (.A(_10201_),
    .Y(_10202_));
 sky130_fd_sc_hd__o22a_2 _24550_ (.A1(_10087_),
    .A2(_10137_),
    .B1(_10078_),
    .B2(_10138_),
    .X(_10203_));
 sky130_fd_sc_hd__a2bb2o_2 _24551_ (.A1_N(_10008_),
    .A2_N(_10203_),
    .B1(_10008_),
    .B2(_10203_),
    .X(_10204_));
 sky130_fd_sc_hd__a2bb2o_2 _24552_ (.A1_N(_10006_),
    .A2_N(_10204_),
    .B1(_10006_),
    .B2(_10204_),
    .X(_10205_));
 sky130_vsdinv _24553_ (.A(_10205_),
    .Y(_10206_));
 sky130_fd_sc_hd__a22o_2 _24554_ (.A1(_10202_),
    .A2(_10205_),
    .B1(_10201_),
    .B2(_10206_),
    .X(_10207_));
 sky130_fd_sc_hd__o22a_2 _24555_ (.A1(_10140_),
    .A2(_10141_),
    .B1(_10143_),
    .B2(_10146_),
    .X(_10208_));
 sky130_fd_sc_hd__a2bb2o_2 _24556_ (.A1_N(_10207_),
    .A2_N(_10208_),
    .B1(_10207_),
    .B2(_10208_),
    .X(_10209_));
 sky130_fd_sc_hd__buf_1 _24557_ (.A(_10028_),
    .X(_10210_));
 sky130_fd_sc_hd__o22a_2 _24558_ (.A1(_10018_),
    .A2(_10144_),
    .B1(_10151_),
    .B2(_10145_),
    .X(_10211_));
 sky130_fd_sc_hd__a2bb2o_2 _24559_ (.A1_N(_10026_),
    .A2_N(_10211_),
    .B1(_10026_),
    .B2(_10211_),
    .X(_10212_));
 sky130_fd_sc_hd__a2bb2o_2 _24560_ (.A1_N(_10210_),
    .A2_N(_10212_),
    .B1(_10016_),
    .B2(_10212_),
    .X(_10213_));
 sky130_fd_sc_hd__a2bb2o_2 _24561_ (.A1_N(_10209_),
    .A2_N(_10213_),
    .B1(_10209_),
    .B2(_10213_),
    .X(_10214_));
 sky130_fd_sc_hd__o22a_2 _24562_ (.A1(_10148_),
    .A2(_10149_),
    .B1(_10150_),
    .B2(_10154_),
    .X(_10215_));
 sky130_fd_sc_hd__a2bb2o_2 _24563_ (.A1_N(_10214_),
    .A2_N(_10215_),
    .B1(_10214_),
    .B2(_10215_),
    .X(_10216_));
 sky130_fd_sc_hd__o22a_2 _24564_ (.A1(_10026_),
    .A2(_10152_),
    .B1(_10028_),
    .B2(_10153_),
    .X(_10217_));
 sky130_fd_sc_hd__or2_2 _24565_ (.A(_09719_),
    .B(_10217_),
    .X(_10218_));
 sky130_fd_sc_hd__a21bo_2 _24566_ (.A1(_10025_),
    .A2(_10217_),
    .B1_N(_10218_),
    .X(_10219_));
 sky130_fd_sc_hd__a2bb2o_2 _24567_ (.A1_N(_10216_),
    .A2_N(_10219_),
    .B1(_10216_),
    .B2(_10219_),
    .X(_10220_));
 sky130_fd_sc_hd__o22a_2 _24568_ (.A1(_10155_),
    .A2(_10156_),
    .B1(_10157_),
    .B2(_10160_),
    .X(_10221_));
 sky130_fd_sc_hd__a2bb2o_2 _24569_ (.A1_N(_10220_),
    .A2_N(_10221_),
    .B1(_10220_),
    .B2(_10221_),
    .X(_10222_));
 sky130_fd_sc_hd__a2bb2o_2 _24570_ (.A1_N(_10159_),
    .A2_N(_10222_),
    .B1(_10159_),
    .B2(_10222_),
    .X(_10223_));
 sky130_fd_sc_hd__o22a_2 _24571_ (.A1(_10161_),
    .A2(_10162_),
    .B1(_10102_),
    .B2(_10163_),
    .X(_10224_));
 sky130_fd_sc_hd__and2_2 _24572_ (.A(_10223_),
    .B(_10224_),
    .X(_10225_));
 sky130_fd_sc_hd__or2_2 _24573_ (.A(_10223_),
    .B(_10224_),
    .X(_10226_));
 sky130_fd_sc_hd__or2b_2 _24574_ (.A(_10225_),
    .B_N(_10226_),
    .X(_10227_));
 sky130_fd_sc_hd__o21ai_2 _24575_ (.A1(_10167_),
    .A2(_10169_),
    .B1(_10166_),
    .Y(_10228_));
 sky130_fd_sc_hd__a2bb2o_2 _24576_ (.A1_N(_10227_),
    .A2_N(_10228_),
    .B1(_10227_),
    .B2(_10228_),
    .X(_02678_));
 sky130_fd_sc_hd__and4_2 _24577_ (.A(_10044_),
    .B(_09902_),
    .C(_11563_),
    .D(_11881_),
    .X(_10229_));
 sky130_fd_sc_hd__o22a_2 _24578_ (.A1(_10600_),
    .A2(_11883_),
    .B1(_10046_),
    .B2(_09972_),
    .X(_10230_));
 sky130_fd_sc_hd__nor2_2 _24579_ (.A(_10229_),
    .B(_10230_),
    .Y(_10231_));
 sky130_fd_sc_hd__nor2_2 _24580_ (.A(_10049_),
    .B(_10057_),
    .Y(_10232_));
 sky130_fd_sc_hd__a2bb2o_2 _24581_ (.A1_N(_10231_),
    .A2_N(_10232_),
    .B1(_10231_),
    .B2(_10232_),
    .X(_10233_));
 sky130_fd_sc_hd__a21oi_2 _24582_ (.A1(_10172_),
    .A2(_10173_),
    .B1(_10170_),
    .Y(_10234_));
 sky130_fd_sc_hd__o2bb2ai_2 _24583_ (.A1_N(_10233_),
    .A2_N(_10234_),
    .B1(_10233_),
    .B2(_10234_),
    .Y(_10235_));
 sky130_fd_sc_hd__buf_1 _24584_ (.A(_10181_),
    .X(_10236_));
 sky130_fd_sc_hd__nor2_2 _24585_ (.A(_09968_),
    .B(_10066_),
    .Y(_10237_));
 sky130_fd_sc_hd__or2_2 _24586_ (.A(_10589_),
    .B(_09898_),
    .X(_10238_));
 sky130_vsdinv _24587_ (.A(_10238_),
    .Y(_10239_));
 sky130_fd_sc_hd__a2bb2o_2 _24588_ (.A1_N(_10237_),
    .A2_N(_10239_),
    .B1(_10237_),
    .B2(_10239_),
    .X(_10240_));
 sky130_fd_sc_hd__a2bb2o_2 _24589_ (.A1_N(_10236_),
    .A2_N(_10240_),
    .B1(_10236_),
    .B2(_10240_),
    .X(_10241_));
 sky130_fd_sc_hd__o2bb2ai_2 _24590_ (.A1_N(_10235_),
    .A2_N(_10241_),
    .B1(_10235_),
    .B2(_10241_),
    .Y(_10242_));
 sky130_fd_sc_hd__o22a_2 _24591_ (.A1(_10174_),
    .A2(_10175_),
    .B1(_10176_),
    .B2(_10182_),
    .X(_10243_));
 sky130_fd_sc_hd__o2bb2ai_2 _24592_ (.A1_N(_10242_),
    .A2_N(_10243_),
    .B1(_10242_),
    .B2(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__buf_1 _24593_ (.A(_10187_),
    .X(_10245_));
 sky130_fd_sc_hd__o21ba_2 _24594_ (.A1(_10179_),
    .A2(_10236_),
    .B1_N(_10178_),
    .X(_10246_));
 sky130_fd_sc_hd__a2bb2o_2 _24595_ (.A1_N(_10195_),
    .A2_N(_10246_),
    .B1(_10195_),
    .B2(_10246_),
    .X(_10247_));
 sky130_fd_sc_hd__a2bb2o_2 _24596_ (.A1_N(_10245_),
    .A2_N(_10247_),
    .B1(_10245_),
    .B2(_10247_),
    .X(_10248_));
 sky130_fd_sc_hd__o2bb2ai_2 _24597_ (.A1_N(_10244_),
    .A2_N(_10248_),
    .B1(_10244_),
    .B2(_10248_),
    .Y(_10249_));
 sky130_fd_sc_hd__o22a_2 _24598_ (.A1(_10183_),
    .A2(_10184_),
    .B1(_10185_),
    .B2(_10190_),
    .X(_10250_));
 sky130_fd_sc_hd__o2bb2ai_2 _24599_ (.A1_N(_10249_),
    .A2_N(_10250_),
    .B1(_10249_),
    .B2(_10250_),
    .Y(_10251_));
 sky130_fd_sc_hd__buf_1 _24600_ (.A(_10195_),
    .X(_10252_));
 sky130_fd_sc_hd__o22a_2 _24601_ (.A1(_10252_),
    .A2(_10188_),
    .B1(_10187_),
    .B2(_10189_),
    .X(_10253_));
 sky130_fd_sc_hd__a2bb2o_2 _24602_ (.A1_N(_10087_),
    .A2_N(_10253_),
    .B1(_10087_),
    .B2(_10253_),
    .X(_10254_));
 sky130_fd_sc_hd__a2bb2o_2 _24603_ (.A1_N(_10194_),
    .A2_N(_10254_),
    .B1(_10194_),
    .B2(_10254_),
    .X(_10255_));
 sky130_fd_sc_hd__o2bb2ai_2 _24604_ (.A1_N(_10251_),
    .A2_N(_10255_),
    .B1(_10251_),
    .B2(_10255_),
    .Y(_10256_));
 sky130_fd_sc_hd__o22a_2 _24605_ (.A1(_10191_),
    .A2(_10192_),
    .B1(_10193_),
    .B2(_10198_),
    .X(_10257_));
 sky130_fd_sc_hd__o2bb2a_2 _24606_ (.A1_N(_10256_),
    .A2_N(_10257_),
    .B1(_10256_),
    .B2(_10257_),
    .X(_10258_));
 sky130_vsdinv _24607_ (.A(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__buf_1 _24608_ (.A(_10151_),
    .X(_10260_));
 sky130_fd_sc_hd__buf_1 _24609_ (.A(_10008_),
    .X(_10261_));
 sky130_fd_sc_hd__buf_1 _24610_ (.A(_10087_),
    .X(_10262_));
 sky130_fd_sc_hd__buf_1 _24611_ (.A(_10194_),
    .X(_10263_));
 sky130_fd_sc_hd__o22a_2 _24612_ (.A1(_10262_),
    .A2(_10196_),
    .B1(_10263_),
    .B2(_10197_),
    .X(_10264_));
 sky130_fd_sc_hd__a2bb2o_2 _24613_ (.A1_N(_10261_),
    .A2_N(_10264_),
    .B1(_10018_),
    .B2(_10264_),
    .X(_10265_));
 sky130_fd_sc_hd__a2bb2o_2 _24614_ (.A1_N(_10260_),
    .A2_N(_10265_),
    .B1(_10151_),
    .B2(_10265_),
    .X(_10266_));
 sky130_vsdinv _24615_ (.A(_10266_),
    .Y(_10267_));
 sky130_fd_sc_hd__a22o_2 _24616_ (.A1(_10259_),
    .A2(_10266_),
    .B1(_10258_),
    .B2(_10267_),
    .X(_10268_));
 sky130_fd_sc_hd__o22a_2 _24617_ (.A1(_10199_),
    .A2(_10200_),
    .B1(_10202_),
    .B2(_10205_),
    .X(_10269_));
 sky130_fd_sc_hd__a2bb2o_2 _24618_ (.A1_N(_10268_),
    .A2_N(_10269_),
    .B1(_10268_),
    .B2(_10269_),
    .X(_10270_));
 sky130_fd_sc_hd__buf_1 _24619_ (.A(_10210_),
    .X(_10271_));
 sky130_fd_sc_hd__o22a_2 _24620_ (.A1(_10261_),
    .A2(_10203_),
    .B1(_10260_),
    .B2(_10204_),
    .X(_10272_));
 sky130_fd_sc_hd__a2bb2o_2 _24621_ (.A1_N(_10027_),
    .A2_N(_10272_),
    .B1(_10027_),
    .B2(_10272_),
    .X(_10273_));
 sky130_fd_sc_hd__a2bb2o_2 _24622_ (.A1_N(_10271_),
    .A2_N(_10273_),
    .B1(_10271_),
    .B2(_10273_),
    .X(_10274_));
 sky130_fd_sc_hd__a2bb2o_2 _24623_ (.A1_N(_10270_),
    .A2_N(_10274_),
    .B1(_10270_),
    .B2(_10274_),
    .X(_10275_));
 sky130_fd_sc_hd__o22a_2 _24624_ (.A1(_10207_),
    .A2(_10208_),
    .B1(_10209_),
    .B2(_10213_),
    .X(_10276_));
 sky130_fd_sc_hd__a2bb2o_2 _24625_ (.A1_N(_10275_),
    .A2_N(_10276_),
    .B1(_10275_),
    .B2(_10276_),
    .X(_10277_));
 sky130_fd_sc_hd__buf_1 _24626_ (.A(_10025_),
    .X(_10278_));
 sky130_fd_sc_hd__buf_1 _24627_ (.A(_10027_),
    .X(_10279_));
 sky130_fd_sc_hd__o22a_2 _24628_ (.A1(_10279_),
    .A2(_10211_),
    .B1(_10271_),
    .B2(_10212_),
    .X(_10280_));
 sky130_fd_sc_hd__or2_2 _24629_ (.A(_10278_),
    .B(_10280_),
    .X(_10281_));
 sky130_fd_sc_hd__a21bo_2 _24630_ (.A1(_10278_),
    .A2(_10280_),
    .B1_N(_10281_),
    .X(_10282_));
 sky130_fd_sc_hd__a2bb2o_2 _24631_ (.A1_N(_10277_),
    .A2_N(_10282_),
    .B1(_10277_),
    .B2(_10282_),
    .X(_10283_));
 sky130_fd_sc_hd__o22a_2 _24632_ (.A1(_10214_),
    .A2(_10215_),
    .B1(_10216_),
    .B2(_10219_),
    .X(_10284_));
 sky130_fd_sc_hd__a2bb2o_2 _24633_ (.A1_N(_10283_),
    .A2_N(_10284_),
    .B1(_10283_),
    .B2(_10284_),
    .X(_10285_));
 sky130_fd_sc_hd__a2bb2o_2 _24634_ (.A1_N(_10218_),
    .A2_N(_10285_),
    .B1(_10218_),
    .B2(_10285_),
    .X(_10286_));
 sky130_fd_sc_hd__o22a_2 _24635_ (.A1(_10220_),
    .A2(_10221_),
    .B1(_10159_),
    .B2(_10222_),
    .X(_10287_));
 sky130_fd_sc_hd__or2_2 _24636_ (.A(_10286_),
    .B(_10287_),
    .X(_10288_));
 sky130_vsdinv _24637_ (.A(_10288_),
    .Y(_10289_));
 sky130_fd_sc_hd__a21oi_2 _24638_ (.A1(_10286_),
    .A2(_10287_),
    .B1(_10289_),
    .Y(_10290_));
 sky130_vsdinv _24639_ (.A(_10290_),
    .Y(_10291_));
 sky130_fd_sc_hd__or2_2 _24640_ (.A(_10167_),
    .B(_10227_),
    .X(_10292_));
 sky130_fd_sc_hd__o221a_2 _24641_ (.A1(_10166_),
    .A2(_10225_),
    .B1(_10168_),
    .B2(_10292_),
    .C1(_10226_),
    .X(_10293_));
 sky130_fd_sc_hd__o41a_2 _24642_ (.A1(_10038_),
    .A2(_10110_),
    .A3(_10292_),
    .A4(_10043_),
    .B1(_10293_),
    .X(_10294_));
 sky130_vsdinv _24643_ (.A(_10294_),
    .Y(_10295_));
 sky130_fd_sc_hd__o22a_2 _24644_ (.A1(_10291_),
    .A2(_10294_),
    .B1(_10290_),
    .B2(_10295_),
    .X(_02679_));
 sky130_fd_sc_hd__and4_2 _24645_ (.A(_10044_),
    .B(_09972_),
    .C(_11563_),
    .D(_11879_),
    .X(_10296_));
 sky130_fd_sc_hd__o22a_2 _24646_ (.A1(_10599_),
    .A2(_11881_),
    .B1(_10046_),
    .B2(_10057_),
    .X(_10297_));
 sky130_fd_sc_hd__nor2_2 _24647_ (.A(_10296_),
    .B(_10297_),
    .Y(_10298_));
 sky130_fd_sc_hd__nor2_2 _24648_ (.A(_10049_),
    .B(_10066_),
    .Y(_10299_));
 sky130_fd_sc_hd__a2bb2o_2 _24649_ (.A1_N(_10298_),
    .A2_N(_10299_),
    .B1(_10298_),
    .B2(_10299_),
    .X(_10300_));
 sky130_fd_sc_hd__a21oi_2 _24650_ (.A1(_10231_),
    .A2(_10232_),
    .B1(_10229_),
    .Y(_10301_));
 sky130_fd_sc_hd__o2bb2ai_2 _24651_ (.A1_N(_10300_),
    .A2_N(_10301_),
    .B1(_10300_),
    .B2(_10301_),
    .Y(_10302_));
 sky130_fd_sc_hd__or2_2 _24652_ (.A(_10589_),
    .B(_09968_),
    .X(_10303_));
 sky130_fd_sc_hd__a32o_2 _24653_ (.A1(_09980_),
    .A2(_11569_),
    .A3(_10239_),
    .B1(_10238_),
    .B2(_10303_),
    .X(_10304_));
 sky130_fd_sc_hd__a2bb2o_2 _24654_ (.A1_N(_10236_),
    .A2_N(_10304_),
    .B1(_10181_),
    .B2(_10304_),
    .X(_10305_));
 sky130_fd_sc_hd__buf_1 _24655_ (.A(_10305_),
    .X(_10306_));
 sky130_fd_sc_hd__o2bb2ai_2 _24656_ (.A1_N(_10302_),
    .A2_N(_10306_),
    .B1(_10302_),
    .B2(_10306_),
    .Y(_10307_));
 sky130_fd_sc_hd__o22a_2 _24657_ (.A1(_10233_),
    .A2(_10234_),
    .B1(_10235_),
    .B2(_10241_),
    .X(_10308_));
 sky130_fd_sc_hd__o2bb2ai_2 _24658_ (.A1_N(_10307_),
    .A2_N(_10308_),
    .B1(_10307_),
    .B2(_10308_),
    .Y(_10309_));
 sky130_fd_sc_hd__o32a_2 _24659_ (.A1(_09968_),
    .A2(_10066_),
    .A3(_10238_),
    .B1(_10236_),
    .B2(_10240_),
    .X(_10310_));
 sky130_fd_sc_hd__a2bb2o_2 _24660_ (.A1_N(_10252_),
    .A2_N(_10310_),
    .B1(_10252_),
    .B2(_10310_),
    .X(_10311_));
 sky130_fd_sc_hd__a2bb2o_2 _24661_ (.A1_N(_10245_),
    .A2_N(_10311_),
    .B1(_10245_),
    .B2(_10311_),
    .X(_10312_));
 sky130_fd_sc_hd__o2bb2ai_2 _24662_ (.A1_N(_10309_),
    .A2_N(_10312_),
    .B1(_10309_),
    .B2(_10312_),
    .Y(_10313_));
 sky130_fd_sc_hd__o22a_2 _24663_ (.A1(_10242_),
    .A2(_10243_),
    .B1(_10244_),
    .B2(_10248_),
    .X(_10314_));
 sky130_fd_sc_hd__o2bb2ai_2 _24664_ (.A1_N(_10313_),
    .A2_N(_10314_),
    .B1(_10313_),
    .B2(_10314_),
    .Y(_10315_));
 sky130_fd_sc_hd__o22a_2 _24665_ (.A1(_10252_),
    .A2(_10246_),
    .B1(_10187_),
    .B2(_10247_),
    .X(_10316_));
 sky130_fd_sc_hd__a2bb2o_2 _24666_ (.A1_N(_10262_),
    .A2_N(_10316_),
    .B1(_10087_),
    .B2(_10316_),
    .X(_10317_));
 sky130_fd_sc_hd__a2bb2o_2 _24667_ (.A1_N(_10263_),
    .A2_N(_10317_),
    .B1(_10263_),
    .B2(_10317_),
    .X(_10318_));
 sky130_fd_sc_hd__o2bb2ai_2 _24668_ (.A1_N(_10315_),
    .A2_N(_10318_),
    .B1(_10315_),
    .B2(_10318_),
    .Y(_10319_));
 sky130_fd_sc_hd__o22a_2 _24669_ (.A1(_10249_),
    .A2(_10250_),
    .B1(_10251_),
    .B2(_10255_),
    .X(_10320_));
 sky130_fd_sc_hd__o2bb2a_2 _24670_ (.A1_N(_10319_),
    .A2_N(_10320_),
    .B1(_10319_),
    .B2(_10320_),
    .X(_10321_));
 sky130_vsdinv _24671_ (.A(_10321_),
    .Y(_10322_));
 sky130_fd_sc_hd__o22a_2 _24672_ (.A1(_10262_),
    .A2(_10253_),
    .B1(_10194_),
    .B2(_10254_),
    .X(_10323_));
 sky130_fd_sc_hd__a2bb2o_2 _24673_ (.A1_N(_10018_),
    .A2_N(_10323_),
    .B1(_10018_),
    .B2(_10323_),
    .X(_10324_));
 sky130_fd_sc_hd__a2bb2o_2 _24674_ (.A1_N(_10151_),
    .A2_N(_10324_),
    .B1(_10151_),
    .B2(_10324_),
    .X(_10325_));
 sky130_vsdinv _24675_ (.A(_10325_),
    .Y(_10326_));
 sky130_fd_sc_hd__a22o_2 _24676_ (.A1(_10322_),
    .A2(_10325_),
    .B1(_10321_),
    .B2(_10326_),
    .X(_10327_));
 sky130_fd_sc_hd__o22a_2 _24677_ (.A1(_10256_),
    .A2(_10257_),
    .B1(_10259_),
    .B2(_10266_),
    .X(_10328_));
 sky130_fd_sc_hd__a2bb2o_2 _24678_ (.A1_N(_10327_),
    .A2_N(_10328_),
    .B1(_10327_),
    .B2(_10328_),
    .X(_10329_));
 sky130_fd_sc_hd__o22a_2 _24679_ (.A1(_10261_),
    .A2(_10264_),
    .B1(_10260_),
    .B2(_10265_),
    .X(_10330_));
 sky130_fd_sc_hd__a2bb2o_2 _24680_ (.A1_N(_10027_),
    .A2_N(_10330_),
    .B1(_10027_),
    .B2(_10330_),
    .X(_10331_));
 sky130_fd_sc_hd__a2bb2o_2 _24681_ (.A1_N(_10271_),
    .A2_N(_10331_),
    .B1(_10210_),
    .B2(_10331_),
    .X(_10332_));
 sky130_fd_sc_hd__a2bb2o_2 _24682_ (.A1_N(_10329_),
    .A2_N(_10332_),
    .B1(_10329_),
    .B2(_10332_),
    .X(_10333_));
 sky130_fd_sc_hd__o22a_2 _24683_ (.A1(_10268_),
    .A2(_10269_),
    .B1(_10270_),
    .B2(_10274_),
    .X(_10334_));
 sky130_fd_sc_hd__a2bb2o_2 _24684_ (.A1_N(_10333_),
    .A2_N(_10334_),
    .B1(_10333_),
    .B2(_10334_),
    .X(_10335_));
 sky130_fd_sc_hd__o22a_2 _24685_ (.A1(_10279_),
    .A2(_10272_),
    .B1(_10210_),
    .B2(_10273_),
    .X(_10336_));
 sky130_fd_sc_hd__or2_2 _24686_ (.A(_10278_),
    .B(_10336_),
    .X(_10337_));
 sky130_fd_sc_hd__a21bo_2 _24687_ (.A1(_10278_),
    .A2(_10336_),
    .B1_N(_10337_),
    .X(_10338_));
 sky130_fd_sc_hd__a2bb2o_2 _24688_ (.A1_N(_10335_),
    .A2_N(_10338_),
    .B1(_10335_),
    .B2(_10338_),
    .X(_10339_));
 sky130_fd_sc_hd__o22a_2 _24689_ (.A1(_10275_),
    .A2(_10276_),
    .B1(_10277_),
    .B2(_10282_),
    .X(_10340_));
 sky130_fd_sc_hd__a2bb2o_2 _24690_ (.A1_N(_10339_),
    .A2_N(_10340_),
    .B1(_10339_),
    .B2(_10340_),
    .X(_10341_));
 sky130_fd_sc_hd__a2bb2o_2 _24691_ (.A1_N(_10281_),
    .A2_N(_10341_),
    .B1(_10281_),
    .B2(_10341_),
    .X(_10342_));
 sky130_fd_sc_hd__o22a_2 _24692_ (.A1(_10283_),
    .A2(_10284_),
    .B1(_10218_),
    .B2(_10285_),
    .X(_10343_));
 sky130_fd_sc_hd__nor2_2 _24693_ (.A(_10342_),
    .B(_10343_),
    .Y(_10344_));
 sky130_fd_sc_hd__a21oi_2 _24694_ (.A1(_10342_),
    .A2(_10343_),
    .B1(_10344_),
    .Y(_10345_));
 sky130_vsdinv _24695_ (.A(_10345_),
    .Y(_10346_));
 sky130_fd_sc_hd__o21ai_2 _24696_ (.A1(_10291_),
    .A2(_10294_),
    .B1(_10288_),
    .Y(_10347_));
 sky130_fd_sc_hd__a2bb2o_2 _24697_ (.A1_N(_10346_),
    .A2_N(_10347_),
    .B1(_10346_),
    .B2(_10347_),
    .X(_02680_));
 sky130_fd_sc_hd__and4_2 _24698_ (.A(_10044_),
    .B(_10057_),
    .C(_11562_),
    .D(_11875_),
    .X(_10348_));
 sky130_fd_sc_hd__o22a_2 _24699_ (.A1(_10599_),
    .A2(_11879_),
    .B1(_09738_),
    .B2(_09699_),
    .X(_10349_));
 sky130_fd_sc_hd__or2_2 _24700_ (.A(_10348_),
    .B(_10349_),
    .X(_10350_));
 sky130_vsdinv _24701_ (.A(_10350_),
    .Y(_10351_));
 sky130_fd_sc_hd__or2_2 _24702_ (.A(_10589_),
    .B(_10049_),
    .X(_10352_));
 sky130_fd_sc_hd__a32o_2 _24703_ (.A1(_09980_),
    .A2(\pcpi_mul.rs2[30] ),
    .A3(_10351_),
    .B1(_10350_),
    .B2(_10352_),
    .X(_10353_));
 sky130_fd_sc_hd__a31o_2 _24704_ (.A1(\pcpi_mul.rs2[30] ),
    .A2(_11875_),
    .A3(_10298_),
    .B1(_10296_),
    .X(_10354_));
 sky130_vsdinv _24705_ (.A(_10354_),
    .Y(_10355_));
 sky130_vsdinv _24706_ (.A(_10353_),
    .Y(_10356_));
 sky130_fd_sc_hd__a22o_2 _24707_ (.A1(_10353_),
    .A2(_10355_),
    .B1(_10356_),
    .B2(_10354_),
    .X(_10357_));
 sky130_fd_sc_hd__a2bb2o_2 _24708_ (.A1_N(_10305_),
    .A2_N(_10357_),
    .B1(_10305_),
    .B2(_10357_),
    .X(_10358_));
 sky130_fd_sc_hd__o22a_2 _24709_ (.A1(_10300_),
    .A2(_10301_),
    .B1(_10302_),
    .B2(_10306_),
    .X(_10359_));
 sky130_fd_sc_hd__o2bb2a_2 _24710_ (.A1_N(_10358_),
    .A2_N(_10359_),
    .B1(_10358_),
    .B2(_10359_),
    .X(_10360_));
 sky130_vsdinv _24711_ (.A(_10360_),
    .Y(_10361_));
 sky130_fd_sc_hd__o22a_2 _24712_ (.A1(_10238_),
    .A2(_10303_),
    .B1(_10236_),
    .B2(_10304_),
    .X(_10362_));
 sky130_fd_sc_hd__a2bb2o_2 _24713_ (.A1_N(_10195_),
    .A2_N(_10362_),
    .B1(_10195_),
    .B2(_10362_),
    .X(_10363_));
 sky130_fd_sc_hd__a2bb2o_2 _24714_ (.A1_N(_10187_),
    .A2_N(_10363_),
    .B1(_10187_),
    .B2(_10363_),
    .X(_10364_));
 sky130_vsdinv _24715_ (.A(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__a22o_2 _24716_ (.A1(_10361_),
    .A2(_10364_),
    .B1(_10360_),
    .B2(_10365_),
    .X(_10366_));
 sky130_fd_sc_hd__o22a_2 _24717_ (.A1(_10307_),
    .A2(_10308_),
    .B1(_10309_),
    .B2(_10312_),
    .X(_10367_));
 sky130_fd_sc_hd__o2bb2ai_2 _24718_ (.A1_N(_10366_),
    .A2_N(_10367_),
    .B1(_10366_),
    .B2(_10367_),
    .Y(_10368_));
 sky130_fd_sc_hd__o22a_2 _24719_ (.A1(_10252_),
    .A2(_10310_),
    .B1(_10245_),
    .B2(_10311_),
    .X(_10369_));
 sky130_fd_sc_hd__a2bb2o_2 _24720_ (.A1_N(_10262_),
    .A2_N(_10369_),
    .B1(_10262_),
    .B2(_10369_),
    .X(_10370_));
 sky130_fd_sc_hd__a2bb2o_2 _24721_ (.A1_N(_10263_),
    .A2_N(_10370_),
    .B1(_10263_),
    .B2(_10370_),
    .X(_10371_));
 sky130_fd_sc_hd__o2bb2ai_2 _24722_ (.A1_N(_10368_),
    .A2_N(_10371_),
    .B1(_10368_),
    .B2(_10371_),
    .Y(_10372_));
 sky130_fd_sc_hd__o22a_2 _24723_ (.A1(_10313_),
    .A2(_10314_),
    .B1(_10315_),
    .B2(_10318_),
    .X(_10373_));
 sky130_fd_sc_hd__o2bb2a_2 _24724_ (.A1_N(_10372_),
    .A2_N(_10373_),
    .B1(_10372_),
    .B2(_10373_),
    .X(_10374_));
 sky130_fd_sc_hd__o22a_2 _24725_ (.A1(_10262_),
    .A2(_10316_),
    .B1(_10263_),
    .B2(_10317_),
    .X(_10375_));
 sky130_fd_sc_hd__a2bb2o_2 _24726_ (.A1_N(_10261_),
    .A2_N(_10375_),
    .B1(_10261_),
    .B2(_10375_),
    .X(_10376_));
 sky130_fd_sc_hd__a2bb2oi_2 _24727_ (.A1_N(_10260_),
    .A2_N(_10376_),
    .B1(_10260_),
    .B2(_10376_),
    .Y(_10377_));
 sky130_fd_sc_hd__a2bb2o_2 _24728_ (.A1_N(_10374_),
    .A2_N(_10377_),
    .B1(_10374_),
    .B2(_10377_),
    .X(_10378_));
 sky130_fd_sc_hd__o22a_2 _24729_ (.A1(_10319_),
    .A2(_10320_),
    .B1(_10322_),
    .B2(_10325_),
    .X(_10379_));
 sky130_fd_sc_hd__a2bb2o_2 _24730_ (.A1_N(_10378_),
    .A2_N(_10379_),
    .B1(_10378_),
    .B2(_10379_),
    .X(_10380_));
 sky130_fd_sc_hd__o22a_2 _24731_ (.A1(_10261_),
    .A2(_10323_),
    .B1(_10260_),
    .B2(_10324_),
    .X(_10381_));
 sky130_fd_sc_hd__a2bb2o_2 _24732_ (.A1_N(_10279_),
    .A2_N(_10381_),
    .B1(_10279_),
    .B2(_10381_),
    .X(_10382_));
 sky130_fd_sc_hd__a2bb2o_2 _24733_ (.A1_N(_10210_),
    .A2_N(_10382_),
    .B1(_10210_),
    .B2(_10382_),
    .X(_10383_));
 sky130_fd_sc_hd__a2bb2o_2 _24734_ (.A1_N(_10380_),
    .A2_N(_10383_),
    .B1(_10380_),
    .B2(_10383_),
    .X(_10384_));
 sky130_fd_sc_hd__o22a_2 _24735_ (.A1(_10327_),
    .A2(_10328_),
    .B1(_10329_),
    .B2(_10332_),
    .X(_10385_));
 sky130_fd_sc_hd__a2bb2o_2 _24736_ (.A1_N(_10384_),
    .A2_N(_10385_),
    .B1(_10384_),
    .B2(_10385_),
    .X(_10386_));
 sky130_fd_sc_hd__o22ai_2 _24737_ (.A1(_10279_),
    .A2(_10330_),
    .B1(_10271_),
    .B2(_10331_),
    .Y(_10387_));
 sky130_fd_sc_hd__or2_2 _24738_ (.A(_10278_),
    .B(_10387_),
    .X(_10388_));
 sky130_fd_sc_hd__a21boi_2 _24739_ (.A1(_10278_),
    .A2(_10387_),
    .B1_N(_10388_),
    .Y(_10389_));
 sky130_fd_sc_hd__a2bb2o_2 _24740_ (.A1_N(_10386_),
    .A2_N(_10389_),
    .B1(_10386_),
    .B2(_10389_),
    .X(_10390_));
 sky130_fd_sc_hd__o22a_2 _24741_ (.A1(_10333_),
    .A2(_10334_),
    .B1(_10335_),
    .B2(_10338_),
    .X(_10391_));
 sky130_fd_sc_hd__a2bb2o_2 _24742_ (.A1_N(_10390_),
    .A2_N(_10391_),
    .B1(_10390_),
    .B2(_10391_),
    .X(_10392_));
 sky130_fd_sc_hd__a2bb2o_2 _24743_ (.A1_N(_10337_),
    .A2_N(_10392_),
    .B1(_10337_),
    .B2(_10392_),
    .X(_10393_));
 sky130_fd_sc_hd__o22a_2 _24744_ (.A1(_10339_),
    .A2(_10340_),
    .B1(_10281_),
    .B2(_10341_),
    .X(_10394_));
 sky130_fd_sc_hd__a2bb2o_2 _24745_ (.A1_N(_10393_),
    .A2_N(_10394_),
    .B1(_10393_),
    .B2(_10394_),
    .X(_10395_));
 sky130_fd_sc_hd__o2bb2a_2 _24746_ (.A1_N(_10342_),
    .A2_N(_10343_),
    .B1(_10289_),
    .B2(_10344_),
    .X(_10396_));
 sky130_fd_sc_hd__a31oi_2 _24747_ (.A1(_10290_),
    .A2(_10345_),
    .A3(_10295_),
    .B1(_10396_),
    .Y(_10397_));
 sky130_fd_sc_hd__a2bb2oi_2 _24748_ (.A1_N(_10395_),
    .A2_N(_10397_),
    .B1(_10395_),
    .B2(_10397_),
    .Y(_02681_));
 sky130_fd_sc_hd__o22a_2 _24749_ (.A1(_10393_),
    .A2(_10394_),
    .B1(_10395_),
    .B2(_10397_),
    .X(_10398_));
 sky130_fd_sc_hd__o22a_2 _24750_ (.A1(_10378_),
    .A2(_10379_),
    .B1(_10380_),
    .B2(_10383_),
    .X(_10399_));
 sky130_fd_sc_hd__o22ai_2 _24751_ (.A1(_10366_),
    .A2(_10367_),
    .B1(_10368_),
    .B2(_10371_),
    .Y(_10400_));
 sky130_fd_sc_hd__o2bb2a_2 _24752_ (.A1_N(_10399_),
    .A2_N(_10400_),
    .B1(_10399_),
    .B2(_10400_),
    .X(_10401_));
 sky130_fd_sc_hd__or2b_2 _24753_ (.A(_09996_),
    .B_N(_10369_),
    .X(_10402_));
 sky130_fd_sc_hd__a2bb2o_2 _24754_ (.A1_N(_09995_),
    .A2_N(_10369_),
    .B1(_09920_),
    .B2(_10402_),
    .X(_10403_));
 sky130_fd_sc_hd__a2bb2o_2 _24755_ (.A1_N(_10306_),
    .A2_N(_10403_),
    .B1(_10306_),
    .B2(_10403_),
    .X(_10404_));
 sky130_vsdinv _24756_ (.A(_10404_),
    .Y(_10405_));
 sky130_fd_sc_hd__a32o_2 _24757_ (.A1(_09980_),
    .A2(\pcpi_mul.rs2[30] ),
    .A3(_10404_),
    .B1(_10352_),
    .B2(_10405_),
    .X(_10406_));
 sky130_vsdinv _24758_ (.A(_10406_),
    .Y(_10407_));
 sky130_fd_sc_hd__a22o_2 _24759_ (.A1(_10365_),
    .A2(_10406_),
    .B1(_10364_),
    .B2(_10407_),
    .X(_10408_));
 sky130_fd_sc_hd__o2bb2a_2 _24760_ (.A1_N(_10401_),
    .A2_N(_10408_),
    .B1(_10401_),
    .B2(_10408_),
    .X(_10409_));
 sky130_fd_sc_hd__o22a_2 _24761_ (.A1(_10252_),
    .A2(_10362_),
    .B1(_10245_),
    .B2(_10363_),
    .X(_10410_));
 sky130_fd_sc_hd__or2_2 _24762_ (.A(_10589_),
    .B(_10046_),
    .X(_10411_));
 sky130_fd_sc_hd__o22a_2 _24763_ (.A1(_09262_),
    .A2(_09377_),
    .B1(_09381_),
    .B2(_09380_),
    .X(_10412_));
 sky130_fd_sc_hd__o22a_2 _24764_ (.A1(_10390_),
    .A2(_10391_),
    .B1(_10337_),
    .B2(_10392_),
    .X(_10413_));
 sky130_fd_sc_hd__o2bb2a_2 _24765_ (.A1_N(_10412_),
    .A2_N(_10413_),
    .B1(_10412_),
    .B2(_10413_),
    .X(_10414_));
 sky130_fd_sc_hd__a2bb2o_2 _24766_ (.A1_N(_10411_),
    .A2_N(_10414_),
    .B1(_10411_),
    .B2(_10414_),
    .X(_10415_));
 sky130_fd_sc_hd__o2bb2a_2 _24767_ (.A1_N(_10410_),
    .A2_N(_10415_),
    .B1(_10410_),
    .B2(_10415_),
    .X(_10416_));
 sky130_fd_sc_hd__o2bb2ai_2 _24768_ (.A1_N(_10409_),
    .A2_N(_10416_),
    .B1(_10409_),
    .B2(_10416_),
    .Y(_10417_));
 sky130_fd_sc_hd__a2bb2o_2 _24769_ (.A1_N(_10372_),
    .A2_N(_10373_),
    .B1(_10374_),
    .B2(_10377_),
    .X(_10418_));
 sky130_fd_sc_hd__o22a_2 _24770_ (.A1(_10358_),
    .A2(_10359_),
    .B1(_10361_),
    .B2(_10364_),
    .X(_10419_));
 sky130_fd_sc_hd__a2bb2oi_2 _24771_ (.A1_N(_10418_),
    .A2_N(_10419_),
    .B1(_10418_),
    .B2(_10419_),
    .Y(_10420_));
 sky130_fd_sc_hd__o2bb2a_2 _24772_ (.A1_N(_10417_),
    .A2_N(_10420_),
    .B1(_10417_),
    .B2(_10420_),
    .X(_10421_));
 sky130_fd_sc_hd__a31o_2 _24773_ (.A1(_09980_),
    .A2(\pcpi_mul.rs2[30] ),
    .A3(_10351_),
    .B1(_10348_),
    .X(_10422_));
 sky130_fd_sc_hd__o22ai_2 _24774_ (.A1(_10384_),
    .A2(_10385_),
    .B1(_10386_),
    .B2(_10389_),
    .Y(_10423_));
 sky130_fd_sc_hd__o22a_2 _24775_ (.A1(_10353_),
    .A2(_10355_),
    .B1(_10306_),
    .B2(_10357_),
    .X(_10424_));
 sky130_fd_sc_hd__or2b_2 _24776_ (.A(_09864_),
    .B_N(_10375_),
    .X(_10425_));
 sky130_fd_sc_hd__a2bb2o_2 _24777_ (.A1_N(_09863_),
    .A2_N(_10375_),
    .B1(_09272_),
    .B2(_10425_),
    .X(_10426_));
 sky130_fd_sc_hd__a2bb2oi_2 _24778_ (.A1_N(_10424_),
    .A2_N(_10426_),
    .B1(_10424_),
    .B2(_10426_),
    .Y(_10427_));
 sky130_fd_sc_hd__a2bb2oi_2 _24779_ (.A1_N(_10423_),
    .A2_N(_10427_),
    .B1(_10423_),
    .B2(_10427_),
    .Y(_10428_));
 sky130_fd_sc_hd__o22a_2 _24780_ (.A1(_10279_),
    .A2(_10381_),
    .B1(_10271_),
    .B2(_10382_),
    .X(_10429_));
 sky130_fd_sc_hd__a2bb2o_2 _24781_ (.A1_N(_10388_),
    .A2_N(_10429_),
    .B1(_10388_),
    .B2(_10429_),
    .X(_10430_));
 sky130_fd_sc_hd__nor2_2 _24782_ (.A(_10600_),
    .B(_11875_),
    .Y(_10431_));
 sky130_fd_sc_hd__o2bb2a_2 _24783_ (.A1_N(_10430_),
    .A2_N(_10431_),
    .B1(_10430_),
    .B2(_10431_),
    .X(_10432_));
 sky130_fd_sc_hd__o2bb2a_2 _24784_ (.A1_N(_10428_),
    .A2_N(_10432_),
    .B1(_10428_),
    .B2(_10432_),
    .X(_10433_));
 sky130_fd_sc_hd__a2bb2o_2 _24785_ (.A1_N(_10422_),
    .A2_N(_10433_),
    .B1(_10422_),
    .B2(_10433_),
    .X(_10434_));
 sky130_fd_sc_hd__nand2_2 _24786_ (.A(_10421_),
    .B(_10434_),
    .Y(_10435_));
 sky130_fd_sc_hd__or2_2 _24787_ (.A(_10421_),
    .B(_10434_),
    .X(_10436_));
 sky130_fd_sc_hd__nand2_2 _24788_ (.A(_10435_),
    .B(_10436_),
    .Y(_10437_));
 sky130_fd_sc_hd__nand2_2 _24789_ (.A(_10398_),
    .B(_10437_),
    .Y(_10438_));
 sky130_fd_sc_hd__or2_2 _24790_ (.A(_10398_),
    .B(_10437_),
    .X(_10439_));
 sky130_fd_sc_hd__and2_2 _24791_ (.A(_10438_),
    .B(_10439_),
    .X(_02682_));
 sky130_fd_sc_hd__or2_2 _24792_ (.A(_04763_),
    .B(_04766_),
    .X(_10440_));
 sky130_fd_sc_hd__a2bb2o_2 _24793_ (.A1_N(_04790_),
    .A2_N(_10440_),
    .B1(_04790_),
    .B2(_10440_),
    .X(_02628_));
 sky130_fd_sc_hd__and2_2 _24794_ (.A(_02318_),
    .B(_00066_),
    .X(_00067_));
 sky130_fd_sc_hd__o21a_2 _24795_ (.A1(instr_sra),
    .A2(instr_srai),
    .B1(_11812_),
    .X(_00216_));
 sky130_fd_sc_hd__o21ai_2 _24796_ (.A1(_10654_),
    .A2(_10646_),
    .B1(_00321_),
    .Y(_10441_));
 sky130_vsdinv _24797_ (.A(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__o221a_2 _24798_ (.A1(_12369_),
    .A2(_10441_),
    .B1(irq_active),
    .B2(_10442_),
    .C1(_11106_),
    .X(_04072_));
 sky130_fd_sc_hd__conb_1 _24799_ (.LO(mem_addr[0]));
 sky130_fd_sc_hd__conb_1 _24800_ (.LO(mem_addr[1]));
 sky130_fd_sc_hd__conb_1 _24801_ (.LO(mem_la_addr[0]));
 sky130_fd_sc_hd__conb_1 _24802_ (.LO(mem_la_addr[1]));
 sky130_fd_sc_hd__conb_1 _24803_ (.LO(trace_data[0]));
 sky130_fd_sc_hd__conb_1 _24804_ (.LO(trace_data[1]));
 sky130_fd_sc_hd__conb_1 _24805_ (.LO(trace_data[2]));
 sky130_fd_sc_hd__conb_1 _24806_ (.LO(trace_data[3]));
 sky130_fd_sc_hd__conb_1 _24807_ (.LO(trace_data[4]));
 sky130_fd_sc_hd__conb_1 _24808_ (.LO(trace_data[5]));
 sky130_fd_sc_hd__conb_1 _24809_ (.LO(trace_data[6]));
 sky130_fd_sc_hd__conb_1 _24810_ (.LO(trace_data[7]));
 sky130_fd_sc_hd__conb_1 _24811_ (.LO(trace_data[8]));
 sky130_fd_sc_hd__conb_1 _24812_ (.LO(trace_data[9]));
 sky130_fd_sc_hd__conb_1 _24813_ (.LO(trace_data[10]));
 sky130_fd_sc_hd__conb_1 _24814_ (.LO(trace_data[11]));
 sky130_fd_sc_hd__conb_1 _24815_ (.LO(trace_data[12]));
 sky130_fd_sc_hd__conb_1 _24816_ (.LO(trace_data[13]));
 sky130_fd_sc_hd__conb_1 _24817_ (.LO(trace_data[14]));
 sky130_fd_sc_hd__conb_1 _24818_ (.LO(trace_data[15]));
 sky130_fd_sc_hd__conb_1 _24819_ (.LO(trace_data[16]));
 sky130_fd_sc_hd__conb_1 _24820_ (.LO(trace_data[17]));
 sky130_fd_sc_hd__conb_1 _24821_ (.LO(trace_data[18]));
 sky130_fd_sc_hd__conb_1 _24822_ (.LO(trace_data[19]));
 sky130_fd_sc_hd__conb_1 _24823_ (.LO(trace_data[20]));
 sky130_fd_sc_hd__conb_1 _24824_ (.LO(trace_data[21]));
 sky130_fd_sc_hd__conb_1 _24825_ (.LO(trace_data[22]));
 sky130_fd_sc_hd__conb_1 _24826_ (.LO(trace_data[23]));
 sky130_fd_sc_hd__conb_1 _24827_ (.LO(trace_data[24]));
 sky130_fd_sc_hd__conb_1 _24828_ (.LO(trace_data[25]));
 sky130_fd_sc_hd__conb_1 _24829_ (.LO(trace_data[26]));
 sky130_fd_sc_hd__conb_1 _24830_ (.LO(trace_data[27]));
 sky130_fd_sc_hd__conb_1 _24831_ (.LO(trace_data[28]));
 sky130_fd_sc_hd__conb_1 _24832_ (.LO(trace_data[29]));
 sky130_fd_sc_hd__conb_1 _24833_ (.LO(trace_data[30]));
 sky130_fd_sc_hd__conb_1 _24834_ (.LO(trace_data[31]));
 sky130_fd_sc_hd__conb_1 _24835_ (.LO(trace_data[32]));
 sky130_fd_sc_hd__conb_1 _24836_ (.LO(trace_data[33]));
 sky130_fd_sc_hd__conb_1 _24837_ (.LO(trace_data[34]));
 sky130_fd_sc_hd__conb_1 _24838_ (.LO(trace_data[35]));
 sky130_fd_sc_hd__conb_1 _24839_ (.LO(trace_valid));
 sky130_fd_sc_hd__conb_1 _24840_ (.LO(_00313_));
 sky130_fd_sc_hd__buf_2 _24841_ (.A(mem_la_wdata[0]),
    .X(pcpi_rs2[0]));
 sky130_fd_sc_hd__buf_2 _24842_ (.A(mem_la_wdata[1]),
    .X(pcpi_rs2[1]));
 sky130_fd_sc_hd__buf_2 _24843_ (.A(mem_la_wdata[2]),
    .X(pcpi_rs2[2]));
 sky130_fd_sc_hd__buf_2 _24844_ (.A(mem_la_wdata[3]),
    .X(pcpi_rs2[3]));
 sky130_fd_sc_hd__buf_2 _24845_ (.A(mem_la_wdata[4]),
    .X(pcpi_rs2[4]));
 sky130_fd_sc_hd__buf_2 _24846_ (.A(mem_la_wdata[5]),
    .X(pcpi_rs2[5]));
 sky130_fd_sc_hd__buf_2 _24847_ (.A(mem_la_wdata[6]),
    .X(pcpi_rs2[6]));
 sky130_fd_sc_hd__buf_2 _24848_ (.A(mem_la_wdata[7]),
    .X(pcpi_rs2[7]));
 sky130_fd_sc_hd__mux2_1 _24849_ (.A0(decoder_trigger),
    .A1(_02410_),
    .S(_00309_),
    .X(_12946_));
 sky130_fd_sc_hd__mux2_1 _24850_ (.A0(\reg_out[2] ),
    .A1(\reg_next_pc[2] ),
    .S(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _24851_ (.A0(_02184_),
    .A1(pcpi_rs1[2]),
    .S(_00301_),
    .X(mem_la_addr[2]));
 sky130_fd_sc_hd__mux2_1 _24852_ (.A0(\reg_out[3] ),
    .A1(\reg_next_pc[3] ),
    .S(_02183_),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_1 _24853_ (.A0(_02185_),
    .A1(pcpi_rs1[3]),
    .S(_00301_),
    .X(mem_la_addr[3]));
 sky130_fd_sc_hd__mux2_1 _24854_ (.A0(\reg_out[4] ),
    .A1(\reg_next_pc[4] ),
    .S(_02183_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _24855_ (.A0(_02186_),
    .A1(pcpi_rs1[4]),
    .S(_00301_),
    .X(mem_la_addr[4]));
 sky130_fd_sc_hd__mux2_1 _24856_ (.A0(\reg_out[5] ),
    .A1(\reg_next_pc[5] ),
    .S(_02183_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_1 _24857_ (.A0(_02187_),
    .A1(pcpi_rs1[5]),
    .S(_00301_),
    .X(mem_la_addr[5]));
 sky130_fd_sc_hd__mux2_1 _24858_ (.A0(\reg_out[6] ),
    .A1(\reg_next_pc[6] ),
    .S(_02183_),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_1 _24859_ (.A0(_02188_),
    .A1(pcpi_rs1[6]),
    .S(_00301_),
    .X(mem_la_addr[6]));
 sky130_fd_sc_hd__mux2_1 _24860_ (.A0(\reg_out[7] ),
    .A1(\reg_next_pc[7] ),
    .S(_02183_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _24861_ (.A0(_02189_),
    .A1(pcpi_rs1[7]),
    .S(_00301_),
    .X(mem_la_addr[7]));
 sky130_fd_sc_hd__mux2_1 _24862_ (.A0(\reg_out[8] ),
    .A1(\reg_next_pc[8] ),
    .S(_02183_),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_1 _24863_ (.A0(_02190_),
    .A1(pcpi_rs1[8]),
    .S(_00301_),
    .X(mem_la_addr[8]));
 sky130_fd_sc_hd__mux2_1 _24864_ (.A0(\reg_out[9] ),
    .A1(\reg_next_pc[9] ),
    .S(_02183_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _24865_ (.A0(_02191_),
    .A1(pcpi_rs1[9]),
    .S(_00301_),
    .X(mem_la_addr[9]));
 sky130_fd_sc_hd__mux2_1 _24866_ (.A0(\reg_out[10] ),
    .A1(\reg_next_pc[10] ),
    .S(_02183_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_1 _24867_ (.A0(_02192_),
    .A1(pcpi_rs1[10]),
    .S(_00301_),
    .X(mem_la_addr[10]));
 sky130_fd_sc_hd__mux2_1 _24868_ (.A0(\reg_out[11] ),
    .A1(\reg_next_pc[11] ),
    .S(_02183_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_1 _24869_ (.A0(_02193_),
    .A1(pcpi_rs1[11]),
    .S(_00301_),
    .X(mem_la_addr[11]));
 sky130_fd_sc_hd__mux2_1 _24870_ (.A0(\reg_out[12] ),
    .A1(\reg_next_pc[12] ),
    .S(_02183_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_1 _24871_ (.A0(_02194_),
    .A1(pcpi_rs1[12]),
    .S(_00301_),
    .X(mem_la_addr[12]));
 sky130_fd_sc_hd__mux2_1 _24872_ (.A0(\reg_out[13] ),
    .A1(\reg_next_pc[13] ),
    .S(_02183_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_1 _24873_ (.A0(_02195_),
    .A1(pcpi_rs1[13]),
    .S(_00301_),
    .X(mem_la_addr[13]));
 sky130_fd_sc_hd__mux2_1 _24874_ (.A0(\reg_out[14] ),
    .A1(\reg_next_pc[14] ),
    .S(_02183_),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_1 _24875_ (.A0(_02196_),
    .A1(pcpi_rs1[14]),
    .S(_00301_),
    .X(mem_la_addr[14]));
 sky130_fd_sc_hd__mux2_1 _24876_ (.A0(\reg_out[15] ),
    .A1(\reg_next_pc[15] ),
    .S(_02183_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_1 _24877_ (.A0(_02197_),
    .A1(pcpi_rs1[15]),
    .S(_00301_),
    .X(mem_la_addr[15]));
 sky130_fd_sc_hd__mux2_1 _24878_ (.A0(\reg_out[16] ),
    .A1(\reg_next_pc[16] ),
    .S(_02183_),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_1 _24879_ (.A0(_02198_),
    .A1(pcpi_rs1[16]),
    .S(_00301_),
    .X(mem_la_addr[16]));
 sky130_fd_sc_hd__mux2_1 _24880_ (.A0(\reg_out[17] ),
    .A1(\reg_next_pc[17] ),
    .S(_02183_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_1 _24881_ (.A0(_02199_),
    .A1(pcpi_rs1[17]),
    .S(_00301_),
    .X(mem_la_addr[17]));
 sky130_fd_sc_hd__mux2_1 _24882_ (.A0(\reg_out[18] ),
    .A1(\reg_next_pc[18] ),
    .S(_02183_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _24883_ (.A0(_02200_),
    .A1(pcpi_rs1[18]),
    .S(_00301_),
    .X(mem_la_addr[18]));
 sky130_fd_sc_hd__mux2_1 _24884_ (.A0(\reg_out[19] ),
    .A1(\reg_next_pc[19] ),
    .S(_02183_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _24885_ (.A0(_02201_),
    .A1(pcpi_rs1[19]),
    .S(_00301_),
    .X(mem_la_addr[19]));
 sky130_fd_sc_hd__mux2_1 _24886_ (.A0(\reg_out[20] ),
    .A1(\reg_next_pc[20] ),
    .S(_02183_),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_1 _24887_ (.A0(_02202_),
    .A1(pcpi_rs1[20]),
    .S(_00301_),
    .X(mem_la_addr[20]));
 sky130_fd_sc_hd__mux2_1 _24888_ (.A0(\reg_out[21] ),
    .A1(\reg_next_pc[21] ),
    .S(_02183_),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_1 _24889_ (.A0(_02203_),
    .A1(pcpi_rs1[21]),
    .S(_00301_),
    .X(mem_la_addr[21]));
 sky130_fd_sc_hd__mux2_1 _24890_ (.A0(\reg_out[22] ),
    .A1(\reg_next_pc[22] ),
    .S(_02183_),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_1 _24891_ (.A0(_02204_),
    .A1(pcpi_rs1[22]),
    .S(_00301_),
    .X(mem_la_addr[22]));
 sky130_fd_sc_hd__mux2_1 _24892_ (.A0(\reg_out[23] ),
    .A1(\reg_next_pc[23] ),
    .S(_02183_),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_1 _24893_ (.A0(_02205_),
    .A1(pcpi_rs1[23]),
    .S(_00301_),
    .X(mem_la_addr[23]));
 sky130_fd_sc_hd__mux2_1 _24894_ (.A0(\reg_out[24] ),
    .A1(\reg_next_pc[24] ),
    .S(_02183_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _24895_ (.A0(_02206_),
    .A1(pcpi_rs1[24]),
    .S(_00301_),
    .X(mem_la_addr[24]));
 sky130_fd_sc_hd__mux2_1 _24896_ (.A0(\reg_out[25] ),
    .A1(\reg_next_pc[25] ),
    .S(_02183_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _24897_ (.A0(_02207_),
    .A1(pcpi_rs1[25]),
    .S(_00301_),
    .X(mem_la_addr[25]));
 sky130_fd_sc_hd__mux2_1 _24898_ (.A0(\reg_out[26] ),
    .A1(\reg_next_pc[26] ),
    .S(_02183_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_1 _24899_ (.A0(_02208_),
    .A1(pcpi_rs1[26]),
    .S(_00301_),
    .X(mem_la_addr[26]));
 sky130_fd_sc_hd__mux2_1 _24900_ (.A0(\reg_out[27] ),
    .A1(\reg_next_pc[27] ),
    .S(_02183_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _24901_ (.A0(_02209_),
    .A1(pcpi_rs1[27]),
    .S(_00301_),
    .X(mem_la_addr[27]));
 sky130_fd_sc_hd__mux2_1 _24902_ (.A0(\reg_out[28] ),
    .A1(\reg_next_pc[28] ),
    .S(_02183_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_1 _24903_ (.A0(_02210_),
    .A1(pcpi_rs1[28]),
    .S(_00301_),
    .X(mem_la_addr[28]));
 sky130_fd_sc_hd__mux2_1 _24904_ (.A0(\reg_out[29] ),
    .A1(\reg_next_pc[29] ),
    .S(_02183_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _24905_ (.A0(_02211_),
    .A1(pcpi_rs1[29]),
    .S(_00301_),
    .X(mem_la_addr[29]));
 sky130_fd_sc_hd__mux2_1 _24906_ (.A0(\reg_out[30] ),
    .A1(\reg_next_pc[30] ),
    .S(_02183_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _24907_ (.A0(_02212_),
    .A1(pcpi_rs1[30]),
    .S(_00301_),
    .X(mem_la_addr[30]));
 sky130_fd_sc_hd__mux2_1 _24908_ (.A0(\reg_out[31] ),
    .A1(\reg_next_pc[31] ),
    .S(_02183_),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_1 _24909_ (.A0(_02213_),
    .A1(pcpi_rs1[31]),
    .S(_00301_),
    .X(mem_la_addr[31]));
 sky130_fd_sc_hd__mux2_1 _24910_ (.A0(_02167_),
    .A1(pcpi_rs2[8]),
    .S(_01683_),
    .X(mem_la_wdata[8]));
 sky130_fd_sc_hd__mux2_1 _24911_ (.A0(_02168_),
    .A1(pcpi_rs2[9]),
    .S(_01683_),
    .X(mem_la_wdata[9]));
 sky130_fd_sc_hd__mux2_1 _24912_ (.A0(_02169_),
    .A1(pcpi_rs2[10]),
    .S(_01683_),
    .X(mem_la_wdata[10]));
 sky130_fd_sc_hd__mux2_1 _24913_ (.A0(_02170_),
    .A1(pcpi_rs2[11]),
    .S(_01683_),
    .X(mem_la_wdata[11]));
 sky130_fd_sc_hd__mux2_1 _24914_ (.A0(_02171_),
    .A1(pcpi_rs2[12]),
    .S(_01683_),
    .X(mem_la_wdata[12]));
 sky130_fd_sc_hd__mux2_1 _24915_ (.A0(_02172_),
    .A1(pcpi_rs2[13]),
    .S(_01683_),
    .X(mem_la_wdata[13]));
 sky130_fd_sc_hd__mux2_1 _24916_ (.A0(_02173_),
    .A1(pcpi_rs2[14]),
    .S(_01683_),
    .X(mem_la_wdata[14]));
 sky130_fd_sc_hd__mux2_1 _24917_ (.A0(_02174_),
    .A1(pcpi_rs2[15]),
    .S(_01683_),
    .X(mem_la_wdata[15]));
 sky130_fd_sc_hd__mux2_1 _24918_ (.A0(_02175_),
    .A1(pcpi_rs2[16]),
    .S(_01683_),
    .X(mem_la_wdata[16]));
 sky130_fd_sc_hd__mux2_1 _24919_ (.A0(_02176_),
    .A1(pcpi_rs2[17]),
    .S(_01683_),
    .X(mem_la_wdata[17]));
 sky130_fd_sc_hd__mux2_1 _24920_ (.A0(_02177_),
    .A1(pcpi_rs2[18]),
    .S(_01683_),
    .X(mem_la_wdata[18]));
 sky130_fd_sc_hd__mux2_1 _24921_ (.A0(_02178_),
    .A1(pcpi_rs2[19]),
    .S(_01683_),
    .X(mem_la_wdata[19]));
 sky130_fd_sc_hd__mux2_1 _24922_ (.A0(_02179_),
    .A1(pcpi_rs2[20]),
    .S(_01683_),
    .X(mem_la_wdata[20]));
 sky130_fd_sc_hd__mux2_1 _24923_ (.A0(_02180_),
    .A1(pcpi_rs2[21]),
    .S(_01683_),
    .X(mem_la_wdata[21]));
 sky130_fd_sc_hd__mux2_1 _24924_ (.A0(_02181_),
    .A1(pcpi_rs2[22]),
    .S(_01683_),
    .X(mem_la_wdata[22]));
 sky130_fd_sc_hd__mux2_1 _24925_ (.A0(_02182_),
    .A1(pcpi_rs2[23]),
    .S(_01683_),
    .X(mem_la_wdata[23]));
 sky130_fd_sc_hd__mux2_1 _24926_ (.A0(_02167_),
    .A1(pcpi_rs2[24]),
    .S(_01683_),
    .X(mem_la_wdata[24]));
 sky130_fd_sc_hd__mux2_1 _24927_ (.A0(_02168_),
    .A1(pcpi_rs2[25]),
    .S(_01683_),
    .X(mem_la_wdata[25]));
 sky130_fd_sc_hd__mux2_1 _24928_ (.A0(_02169_),
    .A1(pcpi_rs2[26]),
    .S(_01683_),
    .X(mem_la_wdata[26]));
 sky130_fd_sc_hd__mux2_1 _24929_ (.A0(_02170_),
    .A1(pcpi_rs2[27]),
    .S(_01683_),
    .X(mem_la_wdata[27]));
 sky130_fd_sc_hd__mux2_1 _24930_ (.A0(_02171_),
    .A1(pcpi_rs2[28]),
    .S(_01683_),
    .X(mem_la_wdata[28]));
 sky130_fd_sc_hd__mux2_1 _24931_ (.A0(_02172_),
    .A1(pcpi_rs2[29]),
    .S(_01683_),
    .X(mem_la_wdata[29]));
 sky130_fd_sc_hd__mux2_1 _24932_ (.A0(_02173_),
    .A1(pcpi_rs2[30]),
    .S(_01683_),
    .X(mem_la_wdata[30]));
 sky130_fd_sc_hd__mux2_1 _24933_ (.A0(_02174_),
    .A1(pcpi_rs2[31]),
    .S(_01683_),
    .X(mem_la_wdata[31]));
 sky130_fd_sc_hd__mux2_1 _24934_ (.A0(\mem_rdata_q[7] ),
    .A1(mem_rdata[7]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[7] ));
 sky130_fd_sc_hd__mux2_1 _24935_ (.A0(\mem_rdata_q[8] ),
    .A1(mem_rdata[8]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[8] ));
 sky130_fd_sc_hd__mux2_1 _24936_ (.A0(\mem_rdata_q[9] ),
    .A1(mem_rdata[9]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[9] ));
 sky130_fd_sc_hd__mux2_1 _24937_ (.A0(\mem_rdata_q[10] ),
    .A1(mem_rdata[10]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[10] ));
 sky130_fd_sc_hd__mux2_1 _24938_ (.A0(\mem_rdata_q[11] ),
    .A1(mem_rdata[11]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[11] ));
 sky130_fd_sc_hd__mux2_1 _24939_ (.A0(\mem_rdata_q[12] ),
    .A1(mem_rdata[12]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[12] ));
 sky130_fd_sc_hd__mux2_1 _24940_ (.A0(\mem_rdata_q[13] ),
    .A1(mem_rdata[13]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[13] ));
 sky130_fd_sc_hd__mux2_1 _24941_ (.A0(\mem_rdata_q[14] ),
    .A1(mem_rdata[14]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[14] ));
 sky130_fd_sc_hd__mux2_1 _24942_ (.A0(\mem_rdata_q[15] ),
    .A1(mem_rdata[15]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[15] ));
 sky130_fd_sc_hd__mux2_1 _24943_ (.A0(\mem_rdata_q[16] ),
    .A1(mem_rdata[16]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[16] ));
 sky130_fd_sc_hd__mux2_1 _24944_ (.A0(\mem_rdata_q[17] ),
    .A1(mem_rdata[17]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[17] ));
 sky130_fd_sc_hd__mux2_1 _24945_ (.A0(\mem_rdata_q[18] ),
    .A1(mem_rdata[18]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[18] ));
 sky130_fd_sc_hd__mux2_1 _24946_ (.A0(\mem_rdata_q[19] ),
    .A1(mem_rdata[19]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[19] ));
 sky130_fd_sc_hd__mux2_1 _24947_ (.A0(\mem_rdata_q[20] ),
    .A1(mem_rdata[20]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[20] ));
 sky130_fd_sc_hd__mux2_1 _24948_ (.A0(\mem_rdata_q[21] ),
    .A1(mem_rdata[21]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[21] ));
 sky130_fd_sc_hd__mux2_1 _24949_ (.A0(\mem_rdata_q[22] ),
    .A1(mem_rdata[22]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[22] ));
 sky130_fd_sc_hd__mux2_1 _24950_ (.A0(\mem_rdata_q[23] ),
    .A1(mem_rdata[23]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[23] ));
 sky130_fd_sc_hd__mux2_1 _24951_ (.A0(\mem_rdata_q[24] ),
    .A1(mem_rdata[24]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[24] ));
 sky130_fd_sc_hd__mux2_1 _24952_ (.A0(\mem_rdata_q[25] ),
    .A1(mem_rdata[25]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[25] ));
 sky130_fd_sc_hd__mux2_1 _24953_ (.A0(\mem_rdata_q[26] ),
    .A1(mem_rdata[26]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[26] ));
 sky130_fd_sc_hd__mux2_1 _24954_ (.A0(\mem_rdata_q[27] ),
    .A1(mem_rdata[27]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[27] ));
 sky130_fd_sc_hd__mux2_1 _24955_ (.A0(\mem_rdata_q[28] ),
    .A1(mem_rdata[28]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[28] ));
 sky130_fd_sc_hd__mux2_1 _24956_ (.A0(\mem_rdata_q[29] ),
    .A1(mem_rdata[29]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[29] ));
 sky130_fd_sc_hd__mux2_1 _24957_ (.A0(\mem_rdata_q[30] ),
    .A1(mem_rdata[30]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[30] ));
 sky130_fd_sc_hd__mux2_1 _24958_ (.A0(\mem_rdata_q[31] ),
    .A1(mem_rdata[31]),
    .S(mem_xfer),
    .X(\mem_rdata_latched[31] ));
 sky130_fd_sc_hd__mux2_1 _24959_ (.A0(_02134_),
    .A1(\alu_add_sub[0] ),
    .S(_02133_),
    .X(\alu_out[0] ));
 sky130_fd_sc_hd__mux2_1 _24960_ (.A0(_02135_),
    .A1(\alu_add_sub[1] ),
    .S(_02133_),
    .X(\alu_out[1] ));
 sky130_fd_sc_hd__mux2_1 _24961_ (.A0(_02136_),
    .A1(\alu_add_sub[2] ),
    .S(_02133_),
    .X(\alu_out[2] ));
 sky130_fd_sc_hd__mux2_1 _24962_ (.A0(_02137_),
    .A1(\alu_add_sub[3] ),
    .S(_02133_),
    .X(\alu_out[3] ));
 sky130_fd_sc_hd__mux2_1 _24963_ (.A0(_02138_),
    .A1(\alu_add_sub[4] ),
    .S(_02133_),
    .X(\alu_out[4] ));
 sky130_fd_sc_hd__mux2_1 _24964_ (.A0(_02139_),
    .A1(\alu_add_sub[5] ),
    .S(_02133_),
    .X(\alu_out[5] ));
 sky130_fd_sc_hd__mux2_1 _24965_ (.A0(_02140_),
    .A1(\alu_add_sub[6] ),
    .S(_02133_),
    .X(\alu_out[6] ));
 sky130_fd_sc_hd__mux2_1 _24966_ (.A0(_02141_),
    .A1(\alu_add_sub[7] ),
    .S(_02133_),
    .X(\alu_out[7] ));
 sky130_fd_sc_hd__mux2_1 _24967_ (.A0(_02142_),
    .A1(\alu_add_sub[8] ),
    .S(_02133_),
    .X(\alu_out[8] ));
 sky130_fd_sc_hd__mux2_1 _24968_ (.A0(_02143_),
    .A1(\alu_add_sub[9] ),
    .S(_02133_),
    .X(\alu_out[9] ));
 sky130_fd_sc_hd__mux2_1 _24969_ (.A0(_02144_),
    .A1(\alu_add_sub[10] ),
    .S(_02133_),
    .X(\alu_out[10] ));
 sky130_fd_sc_hd__mux2_1 _24970_ (.A0(_02145_),
    .A1(\alu_add_sub[11] ),
    .S(_02133_),
    .X(\alu_out[11] ));
 sky130_fd_sc_hd__mux2_1 _24971_ (.A0(_02146_),
    .A1(\alu_add_sub[12] ),
    .S(_02133_),
    .X(\alu_out[12] ));
 sky130_fd_sc_hd__mux2_1 _24972_ (.A0(_02147_),
    .A1(\alu_add_sub[13] ),
    .S(_02133_),
    .X(\alu_out[13] ));
 sky130_fd_sc_hd__mux2_1 _24973_ (.A0(_02148_),
    .A1(\alu_add_sub[14] ),
    .S(_02133_),
    .X(\alu_out[14] ));
 sky130_fd_sc_hd__mux2_1 _24974_ (.A0(_02149_),
    .A1(\alu_add_sub[15] ),
    .S(_02133_),
    .X(\alu_out[15] ));
 sky130_fd_sc_hd__mux2_1 _24975_ (.A0(_02150_),
    .A1(\alu_add_sub[16] ),
    .S(_02133_),
    .X(\alu_out[16] ));
 sky130_fd_sc_hd__mux2_1 _24976_ (.A0(_02151_),
    .A1(\alu_add_sub[17] ),
    .S(_02133_),
    .X(\alu_out[17] ));
 sky130_fd_sc_hd__mux2_1 _24977_ (.A0(_02152_),
    .A1(\alu_add_sub[18] ),
    .S(_02133_),
    .X(\alu_out[18] ));
 sky130_fd_sc_hd__mux2_1 _24978_ (.A0(_02153_),
    .A1(\alu_add_sub[19] ),
    .S(_02133_),
    .X(\alu_out[19] ));
 sky130_fd_sc_hd__mux2_1 _24979_ (.A0(_02154_),
    .A1(\alu_add_sub[20] ),
    .S(_02133_),
    .X(\alu_out[20] ));
 sky130_fd_sc_hd__mux2_1 _24980_ (.A0(_02155_),
    .A1(\alu_add_sub[21] ),
    .S(_02133_),
    .X(\alu_out[21] ));
 sky130_fd_sc_hd__mux2_1 _24981_ (.A0(_02156_),
    .A1(\alu_add_sub[22] ),
    .S(_02133_),
    .X(\alu_out[22] ));
 sky130_fd_sc_hd__mux2_1 _24982_ (.A0(_02157_),
    .A1(\alu_add_sub[23] ),
    .S(_02133_),
    .X(\alu_out[23] ));
 sky130_fd_sc_hd__mux2_1 _24983_ (.A0(_02158_),
    .A1(\alu_add_sub[24] ),
    .S(_02133_),
    .X(\alu_out[24] ));
 sky130_fd_sc_hd__mux2_1 _24984_ (.A0(_02159_),
    .A1(\alu_add_sub[25] ),
    .S(_02133_),
    .X(\alu_out[25] ));
 sky130_fd_sc_hd__mux2_1 _24985_ (.A0(_02160_),
    .A1(\alu_add_sub[26] ),
    .S(_02133_),
    .X(\alu_out[26] ));
 sky130_fd_sc_hd__mux2_1 _24986_ (.A0(_02161_),
    .A1(\alu_add_sub[27] ),
    .S(_02133_),
    .X(\alu_out[27] ));
 sky130_fd_sc_hd__mux2_1 _24987_ (.A0(_02162_),
    .A1(\alu_add_sub[28] ),
    .S(_02133_),
    .X(\alu_out[28] ));
 sky130_fd_sc_hd__mux2_1 _24988_ (.A0(_02163_),
    .A1(\alu_add_sub[29] ),
    .S(_02133_),
    .X(\alu_out[29] ));
 sky130_fd_sc_hd__mux2_1 _24989_ (.A0(_02164_),
    .A1(\alu_add_sub[30] ),
    .S(_02133_),
    .X(\alu_out[30] ));
 sky130_fd_sc_hd__mux2_1 _24990_ (.A0(_02165_),
    .A1(\alu_add_sub[31] ),
    .S(_02133_),
    .X(\alu_out[31] ));
 sky130_fd_sc_hd__mux2_1 _24991_ (.A0(_02071_),
    .A1(\reg_next_pc[0] ),
    .S(_02069_),
    .X(\cpuregs_wrdata[0] ));
 sky130_fd_sc_hd__mux2_1 _24992_ (.A0(_02072_),
    .A1(\reg_pc[1] ),
    .S(_02069_),
    .X(\cpuregs_wrdata[1] ));
 sky130_fd_sc_hd__mux2_1 _24993_ (.A0(_02074_),
    .A1(_02073_),
    .S(_02069_),
    .X(\cpuregs_wrdata[2] ));
 sky130_fd_sc_hd__mux2_1 _24994_ (.A0(_02076_),
    .A1(_02075_),
    .S(_02069_),
    .X(\cpuregs_wrdata[3] ));
 sky130_fd_sc_hd__mux2_1 _24995_ (.A0(_02078_),
    .A1(_02077_),
    .S(_02069_),
    .X(\cpuregs_wrdata[4] ));
 sky130_fd_sc_hd__mux2_1 _24996_ (.A0(_02080_),
    .A1(_02079_),
    .S(_02069_),
    .X(\cpuregs_wrdata[5] ));
 sky130_fd_sc_hd__mux2_1 _24997_ (.A0(_02082_),
    .A1(_02081_),
    .S(_02069_),
    .X(\cpuregs_wrdata[6] ));
 sky130_fd_sc_hd__mux2_1 _24998_ (.A0(_02084_),
    .A1(_02083_),
    .S(_02069_),
    .X(\cpuregs_wrdata[7] ));
 sky130_fd_sc_hd__mux2_1 _24999_ (.A0(_02086_),
    .A1(_02085_),
    .S(_02069_),
    .X(\cpuregs_wrdata[8] ));
 sky130_fd_sc_hd__mux2_1 _25000_ (.A0(_02088_),
    .A1(_02087_),
    .S(_02069_),
    .X(\cpuregs_wrdata[9] ));
 sky130_fd_sc_hd__mux2_1 _25001_ (.A0(_02090_),
    .A1(_02089_),
    .S(_02069_),
    .X(\cpuregs_wrdata[10] ));
 sky130_fd_sc_hd__mux2_1 _25002_ (.A0(_02092_),
    .A1(_02091_),
    .S(_02069_),
    .X(\cpuregs_wrdata[11] ));
 sky130_fd_sc_hd__mux2_1 _25003_ (.A0(_02094_),
    .A1(_02093_),
    .S(_02069_),
    .X(\cpuregs_wrdata[12] ));
 sky130_fd_sc_hd__mux2_1 _25004_ (.A0(_02096_),
    .A1(_02095_),
    .S(_02069_),
    .X(\cpuregs_wrdata[13] ));
 sky130_fd_sc_hd__mux2_1 _25005_ (.A0(_02098_),
    .A1(_02097_),
    .S(_02069_),
    .X(\cpuregs_wrdata[14] ));
 sky130_fd_sc_hd__mux2_1 _25006_ (.A0(_02100_),
    .A1(_02099_),
    .S(_02069_),
    .X(\cpuregs_wrdata[15] ));
 sky130_fd_sc_hd__mux2_1 _25007_ (.A0(_02102_),
    .A1(_02101_),
    .S(_02069_),
    .X(\cpuregs_wrdata[16] ));
 sky130_fd_sc_hd__mux2_1 _25008_ (.A0(_02104_),
    .A1(_02103_),
    .S(_02069_),
    .X(\cpuregs_wrdata[17] ));
 sky130_fd_sc_hd__mux2_1 _25009_ (.A0(_02106_),
    .A1(_02105_),
    .S(_02069_),
    .X(\cpuregs_wrdata[18] ));
 sky130_fd_sc_hd__mux2_1 _25010_ (.A0(_02108_),
    .A1(_02107_),
    .S(_02069_),
    .X(\cpuregs_wrdata[19] ));
 sky130_fd_sc_hd__mux2_1 _25011_ (.A0(_02110_),
    .A1(_02109_),
    .S(_02069_),
    .X(\cpuregs_wrdata[20] ));
 sky130_fd_sc_hd__mux2_1 _25012_ (.A0(_02112_),
    .A1(_02111_),
    .S(_02069_),
    .X(\cpuregs_wrdata[21] ));
 sky130_fd_sc_hd__mux2_1 _25013_ (.A0(_02114_),
    .A1(_02113_),
    .S(_02069_),
    .X(\cpuregs_wrdata[22] ));
 sky130_fd_sc_hd__mux2_1 _25014_ (.A0(_02116_),
    .A1(_02115_),
    .S(_02069_),
    .X(\cpuregs_wrdata[23] ));
 sky130_fd_sc_hd__mux2_1 _25015_ (.A0(_02118_),
    .A1(_02117_),
    .S(_02069_),
    .X(\cpuregs_wrdata[24] ));
 sky130_fd_sc_hd__mux2_1 _25016_ (.A0(_02120_),
    .A1(_02119_),
    .S(_02069_),
    .X(\cpuregs_wrdata[25] ));
 sky130_fd_sc_hd__mux2_1 _25017_ (.A0(_02122_),
    .A1(_02121_),
    .S(_02069_),
    .X(\cpuregs_wrdata[26] ));
 sky130_fd_sc_hd__mux2_1 _25018_ (.A0(_02124_),
    .A1(_02123_),
    .S(_02069_),
    .X(\cpuregs_wrdata[27] ));
 sky130_fd_sc_hd__mux2_1 _25019_ (.A0(_02126_),
    .A1(_02125_),
    .S(_02069_),
    .X(\cpuregs_wrdata[28] ));
 sky130_fd_sc_hd__mux2_1 _25020_ (.A0(_02128_),
    .A1(_02127_),
    .S(_02069_),
    .X(\cpuregs_wrdata[29] ));
 sky130_fd_sc_hd__mux2_1 _25021_ (.A0(_02130_),
    .A1(_02129_),
    .S(_02069_),
    .X(\cpuregs_wrdata[30] ));
 sky130_fd_sc_hd__mux2_1 _25022_ (.A0(_02132_),
    .A1(_02131_),
    .S(_02069_),
    .X(\cpuregs_wrdata[31] ));
 sky130_fd_sc_hd__mux2_1 _25023_ (.A0(_02316_),
    .A1(_02317_),
    .S(_00307_),
    .X(_00004_));
 sky130_fd_sc_hd__mux2_1 _25024_ (.A0(_00347_),
    .A1(_12947_),
    .S(_00336_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _25025_ (.A0(_12947_),
    .A1(_00348_),
    .S(resetn),
    .X(_00003_));
 sky130_fd_sc_hd__mux2_1 _25026_ (.A0(_02304_),
    .A1(_02305_),
    .S(\irq_state[1] ),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _25027_ (.A0(_02306_),
    .A1(_02304_),
    .S(_02217_),
    .X(_00008_));
 sky130_fd_sc_hd__mux2_1 _25028_ (.A0(_02214_),
    .A1(_02215_),
    .S(\irq_state[1] ),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _25029_ (.A0(_02216_),
    .A1(_02214_),
    .S(_02217_),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _25030_ (.A0(_02218_),
    .A1(_02219_),
    .S(\irq_state[1] ),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _25031_ (.A0(_02220_),
    .A1(_02218_),
    .S(_02217_),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _25032_ (.A0(_02221_),
    .A1(_02222_),
    .S(\irq_state[1] ),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _25033_ (.A0(_02223_),
    .A1(_02221_),
    .S(_02217_),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _25034_ (.A0(_02224_),
    .A1(_02225_),
    .S(\irq_state[1] ),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _25035_ (.A0(_02226_),
    .A1(_02224_),
    .S(_02217_),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _25036_ (.A0(_02227_),
    .A1(_02228_),
    .S(\irq_state[1] ),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _25037_ (.A0(_02229_),
    .A1(_02227_),
    .S(_02217_),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _25038_ (.A0(_02230_),
    .A1(_02231_),
    .S(\irq_state[1] ),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _25039_ (.A0(_02232_),
    .A1(_02230_),
    .S(_02217_),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _25040_ (.A0(_02233_),
    .A1(_02234_),
    .S(\irq_state[1] ),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _25041_ (.A0(_02235_),
    .A1(_02233_),
    .S(_02217_),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _25042_ (.A0(_02236_),
    .A1(_02237_),
    .S(\irq_state[1] ),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _25043_ (.A0(_02238_),
    .A1(_02236_),
    .S(_02217_),
    .X(_00009_));
 sky130_fd_sc_hd__mux2_1 _25044_ (.A0(_02239_),
    .A1(_02240_),
    .S(\irq_state[1] ),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _25045_ (.A0(_02241_),
    .A1(_02239_),
    .S(_02217_),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _25046_ (.A0(_02242_),
    .A1(_02243_),
    .S(\irq_state[1] ),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _25047_ (.A0(_02244_),
    .A1(_02242_),
    .S(_02217_),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _25048_ (.A0(_02245_),
    .A1(_02246_),
    .S(\irq_state[1] ),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _25049_ (.A0(_02247_),
    .A1(_02245_),
    .S(_02217_),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _25050_ (.A0(_02248_),
    .A1(_02249_),
    .S(\irq_state[1] ),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _25051_ (.A0(_02250_),
    .A1(_02248_),
    .S(_02217_),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _25052_ (.A0(_02251_),
    .A1(_02252_),
    .S(\irq_state[1] ),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _25053_ (.A0(_02253_),
    .A1(_02251_),
    .S(_02217_),
    .X(_00014_));
 sky130_fd_sc_hd__mux2_1 _25054_ (.A0(_02254_),
    .A1(_02255_),
    .S(\irq_state[1] ),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _25055_ (.A0(_02256_),
    .A1(_02254_),
    .S(_02217_),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _25056_ (.A0(_02257_),
    .A1(_02258_),
    .S(\irq_state[1] ),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _25057_ (.A0(_02259_),
    .A1(_02257_),
    .S(_02217_),
    .X(_00016_));
 sky130_fd_sc_hd__mux2_1 _25058_ (.A0(_02260_),
    .A1(_02261_),
    .S(\irq_state[1] ),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _25059_ (.A0(_02262_),
    .A1(_02260_),
    .S(_02217_),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _25060_ (.A0(_02263_),
    .A1(_02264_),
    .S(\irq_state[1] ),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _25061_ (.A0(_02265_),
    .A1(_02263_),
    .S(_02217_),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _25062_ (.A0(_02266_),
    .A1(_02267_),
    .S(\irq_state[1] ),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _25063_ (.A0(_02268_),
    .A1(_02266_),
    .S(_02217_),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _25064_ (.A0(_02269_),
    .A1(_02270_),
    .S(\irq_state[1] ),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _25065_ (.A0(_02271_),
    .A1(_02269_),
    .S(_02217_),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _25066_ (.A0(_02272_),
    .A1(_02273_),
    .S(\irq_state[1] ),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _25067_ (.A0(_02274_),
    .A1(_02272_),
    .S(_02217_),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _25068_ (.A0(_02275_),
    .A1(_02276_),
    .S(\irq_state[1] ),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _25069_ (.A0(_02277_),
    .A1(_02275_),
    .S(_02217_),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _25070_ (.A0(_02278_),
    .A1(_02279_),
    .S(\irq_state[1] ),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _25071_ (.A0(_02280_),
    .A1(_02278_),
    .S(_02217_),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _25072_ (.A0(_02281_),
    .A1(_02282_),
    .S(\irq_state[1] ),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _25073_ (.A0(_02283_),
    .A1(_02281_),
    .S(_02217_),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _25074_ (.A0(_02284_),
    .A1(_02285_),
    .S(\irq_state[1] ),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _25075_ (.A0(_02286_),
    .A1(_02284_),
    .S(_02217_),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _25076_ (.A0(_02287_),
    .A1(_02288_),
    .S(\irq_state[1] ),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _25077_ (.A0(_02289_),
    .A1(_02287_),
    .S(_02217_),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _25078_ (.A0(_02290_),
    .A1(_02291_),
    .S(\irq_state[1] ),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _25079_ (.A0(_02292_),
    .A1(_02290_),
    .S(_02217_),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _25080_ (.A0(_02293_),
    .A1(_02294_),
    .S(\irq_state[1] ),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _25081_ (.A0(_02295_),
    .A1(_02293_),
    .S(_02217_),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _25082_ (.A0(_02296_),
    .A1(_02297_),
    .S(\irq_state[1] ),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _25083_ (.A0(_02298_),
    .A1(_02296_),
    .S(_02217_),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _25084_ (.A0(_02299_),
    .A1(_02300_),
    .S(\irq_state[1] ),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _25085_ (.A0(_02301_),
    .A1(_02299_),
    .S(_02217_),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_1 _25086_ (.A0(_01467_),
    .A1(\reg_next_pc[1] ),
    .S(_00292_),
    .X(_02590_));
 sky130_fd_sc_hd__mux2_1 _25087_ (.A0(_00295_),
    .A1(\reg_next_pc[2] ),
    .S(_00292_),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_1 _25088_ (.A0(_01470_),
    .A1(\reg_next_pc[3] ),
    .S(_00292_),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_1 _25089_ (.A0(_01478_),
    .A1(\reg_next_pc[5] ),
    .S(_00292_),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_1 _25090_ (.A0(_01481_),
    .A1(\reg_next_pc[6] ),
    .S(_00292_),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_1 _25091_ (.A0(_01484_),
    .A1(\reg_next_pc[7] ),
    .S(_00292_),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_1 _25092_ (.A0(_01487_),
    .A1(\reg_next_pc[8] ),
    .S(_00292_),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_1 _25093_ (.A0(_01490_),
    .A1(\reg_next_pc[9] ),
    .S(_00292_),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_1 _25094_ (.A0(_01493_),
    .A1(\reg_next_pc[10] ),
    .S(_00292_),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_1 _25095_ (.A0(_01496_),
    .A1(\reg_next_pc[11] ),
    .S(_00292_),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_1 _25096_ (.A0(_01499_),
    .A1(\reg_next_pc[12] ),
    .S(_00292_),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_1 _25097_ (.A0(_01502_),
    .A1(\reg_next_pc[13] ),
    .S(_00292_),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_1 _25098_ (.A0(_01505_),
    .A1(\reg_next_pc[14] ),
    .S(_00292_),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_1 _25099_ (.A0(_01508_),
    .A1(\reg_next_pc[15] ),
    .S(_00292_),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_1 _25100_ (.A0(_01511_),
    .A1(\reg_next_pc[16] ),
    .S(_00292_),
    .X(_02565_));
 sky130_fd_sc_hd__mux2_1 _25101_ (.A0(_01514_),
    .A1(\reg_next_pc[17] ),
    .S(_00292_),
    .X(_02566_));
 sky130_fd_sc_hd__mux2_1 _25102_ (.A0(_01517_),
    .A1(\reg_next_pc[18] ),
    .S(_00292_),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_1 _25103_ (.A0(_01520_),
    .A1(\reg_next_pc[19] ),
    .S(_00292_),
    .X(_02568_));
 sky130_fd_sc_hd__mux2_1 _25104_ (.A0(_01523_),
    .A1(\reg_next_pc[20] ),
    .S(_00292_),
    .X(_02569_));
 sky130_fd_sc_hd__mux2_1 _25105_ (.A0(_01526_),
    .A1(\reg_next_pc[21] ),
    .S(_00292_),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_1 _25106_ (.A0(_01529_),
    .A1(\reg_next_pc[22] ),
    .S(_00292_),
    .X(_02572_));
 sky130_fd_sc_hd__mux2_1 _25107_ (.A0(_01532_),
    .A1(\reg_next_pc[23] ),
    .S(_00292_),
    .X(_02573_));
 sky130_fd_sc_hd__mux2_1 _25108_ (.A0(_01535_),
    .A1(\reg_next_pc[24] ),
    .S(_00292_),
    .X(_02574_));
 sky130_fd_sc_hd__mux2_1 _25109_ (.A0(_01538_),
    .A1(\reg_next_pc[25] ),
    .S(_00292_),
    .X(_02575_));
 sky130_fd_sc_hd__mux2_1 _25110_ (.A0(_01541_),
    .A1(\reg_next_pc[26] ),
    .S(_00292_),
    .X(_02576_));
 sky130_fd_sc_hd__mux2_1 _25111_ (.A0(_01544_),
    .A1(\reg_next_pc[27] ),
    .S(_00292_),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_1 _25112_ (.A0(_01547_),
    .A1(\reg_next_pc[28] ),
    .S(_00292_),
    .X(_02578_));
 sky130_fd_sc_hd__mux2_1 _25113_ (.A0(_01550_),
    .A1(\reg_next_pc[29] ),
    .S(_00292_),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_1 _25114_ (.A0(_01553_),
    .A1(\reg_next_pc[30] ),
    .S(_00292_),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_1 _25115_ (.A0(_01556_),
    .A1(\reg_next_pc[31] ),
    .S(_00292_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _25116_ (.A0(_00057_),
    .A1(_00064_),
    .S(mem_la_wdata[3]),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _25117_ (.A0(_00065_),
    .A1(_02543_),
    .S(mem_la_wdata[4]),
    .X(_12983_));
 sky130_fd_sc_hd__mux2_1 _25118_ (.A0(_00075_),
    .A1(_00082_),
    .S(mem_la_wdata[3]),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _25119_ (.A0(_00083_),
    .A1(_02544_),
    .S(mem_la_wdata[4]),
    .X(_12984_));
 sky130_fd_sc_hd__mux2_1 _25120_ (.A0(_00089_),
    .A1(_00092_),
    .S(mem_la_wdata[3]),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _25121_ (.A0(_00093_),
    .A1(_02545_),
    .S(mem_la_wdata[4]),
    .X(_12985_));
 sky130_fd_sc_hd__mux2_1 _25122_ (.A0(_00099_),
    .A1(_00102_),
    .S(mem_la_wdata[3]),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _25123_ (.A0(_00103_),
    .A1(_02546_),
    .S(mem_la_wdata[4]),
    .X(_12986_));
 sky130_fd_sc_hd__mux2_1 _25124_ (.A0(_00107_),
    .A1(_00108_),
    .S(mem_la_wdata[3]),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _25125_ (.A0(_00109_),
    .A1(_02547_),
    .S(mem_la_wdata[4]),
    .X(_12987_));
 sky130_fd_sc_hd__mux2_1 _25126_ (.A0(_00113_),
    .A1(_00114_),
    .S(mem_la_wdata[3]),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _25127_ (.A0(_00115_),
    .A1(_02548_),
    .S(mem_la_wdata[4]),
    .X(_12988_));
 sky130_fd_sc_hd__mux2_1 _25128_ (.A0(_00119_),
    .A1(_00120_),
    .S(mem_la_wdata[3]),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _25129_ (.A0(_00121_),
    .A1(_02549_),
    .S(mem_la_wdata[4]),
    .X(_12989_));
 sky130_fd_sc_hd__mux2_1 _25130_ (.A0(_00125_),
    .A1(_00126_),
    .S(mem_la_wdata[3]),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _25131_ (.A0(_00127_),
    .A1(_02550_),
    .S(mem_la_wdata[4]),
    .X(_12990_));
 sky130_fd_sc_hd__mux2_1 _25132_ (.A0(_00129_),
    .A1(_00106_),
    .S(mem_la_wdata[2]),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _25133_ (.A0(_00130_),
    .A1(_00057_),
    .S(mem_la_wdata[3]),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _25134_ (.A0(_00131_),
    .A1(_02551_),
    .S(mem_la_wdata[4]),
    .X(_12991_));
 sky130_fd_sc_hd__mux2_1 _25135_ (.A0(_00133_),
    .A1(_00112_),
    .S(mem_la_wdata[2]),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _25136_ (.A0(_00134_),
    .A1(_00075_),
    .S(mem_la_wdata[3]),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _25137_ (.A0(_00135_),
    .A1(_02552_),
    .S(mem_la_wdata[4]),
    .X(_12992_));
 sky130_fd_sc_hd__mux2_1 _25138_ (.A0(_00137_),
    .A1(_00118_),
    .S(mem_la_wdata[2]),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _25139_ (.A0(_00138_),
    .A1(_00089_),
    .S(mem_la_wdata[3]),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _25140_ (.A0(_00139_),
    .A1(_02553_),
    .S(mem_la_wdata[4]),
    .X(_12993_));
 sky130_fd_sc_hd__mux2_1 _25141_ (.A0(_00141_),
    .A1(_00124_),
    .S(mem_la_wdata[2]),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _25142_ (.A0(_00142_),
    .A1(_00099_),
    .S(mem_la_wdata[3]),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _25143_ (.A0(_00143_),
    .A1(_02554_),
    .S(mem_la_wdata[4]),
    .X(_12994_));
 sky130_fd_sc_hd__mux2_1 _25144_ (.A0(_00144_),
    .A1(_00136_),
    .S(mem_la_wdata[1]),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _25145_ (.A0(_00145_),
    .A1(_00129_),
    .S(mem_la_wdata[2]),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _25146_ (.A0(_00146_),
    .A1(_00107_),
    .S(mem_la_wdata[3]),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _25147_ (.A0(_00147_),
    .A1(_02555_),
    .S(mem_la_wdata[4]),
    .X(_12995_));
 sky130_fd_sc_hd__mux2_1 _25148_ (.A0(_00148_),
    .A1(_00140_),
    .S(mem_la_wdata[1]),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _25149_ (.A0(_00149_),
    .A1(_00133_),
    .S(mem_la_wdata[2]),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _25150_ (.A0(_00150_),
    .A1(_00113_),
    .S(mem_la_wdata[3]),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _25151_ (.A0(_00151_),
    .A1(_02556_),
    .S(mem_la_wdata[4]),
    .X(_12996_));
 sky130_fd_sc_hd__mux2_1 _25152_ (.A0(pcpi_rs1[30]),
    .A1(pcpi_rs1[29]),
    .S(mem_la_wdata[0]),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _25153_ (.A0(_00152_),
    .A1(_00144_),
    .S(mem_la_wdata[1]),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _25154_ (.A0(_00153_),
    .A1(_00137_),
    .S(mem_la_wdata[2]),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _25155_ (.A0(_00154_),
    .A1(_00119_),
    .S(mem_la_wdata[3]),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _25156_ (.A0(_00155_),
    .A1(_02557_),
    .S(mem_la_wdata[4]),
    .X(_12997_));
 sky130_fd_sc_hd__mux2_1 _25157_ (.A0(pcpi_rs1[31]),
    .A1(pcpi_rs1[30]),
    .S(mem_la_wdata[0]),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _25158_ (.A0(_00156_),
    .A1(_00148_),
    .S(mem_la_wdata[1]),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _25159_ (.A0(_00157_),
    .A1(_00141_),
    .S(mem_la_wdata[2]),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _25160_ (.A0(_00158_),
    .A1(_00125_),
    .S(mem_la_wdata[3]),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _25161_ (.A0(_00159_),
    .A1(_02558_),
    .S(mem_la_wdata[4]),
    .X(_12998_));
 sky130_fd_sc_hd__mux2_1 _25162_ (.A0(pcpi_rs1[0]),
    .A1(pcpi_rs1[1]),
    .S(mem_la_wdata[0]),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _25163_ (.A0(_00160_),
    .A1(_00161_),
    .S(mem_la_wdata[1]),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _25164_ (.A0(_00162_),
    .A1(_00165_),
    .S(mem_la_wdata[2]),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _25165_ (.A0(_00166_),
    .A1(_00173_),
    .S(mem_la_wdata[3]),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _25166_ (.A0(_00174_),
    .A1(_00189_),
    .S(mem_la_wdata[4]),
    .X(_12999_));
 sky130_fd_sc_hd__mux2_1 _25167_ (.A0(pcpi_rs1[1]),
    .A1(pcpi_rs1[2]),
    .S(mem_la_wdata[0]),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _25168_ (.A0(_00190_),
    .A1(_00191_),
    .S(mem_la_wdata[1]),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _25169_ (.A0(_00192_),
    .A1(_00195_),
    .S(mem_la_wdata[2]),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _25170_ (.A0(_00196_),
    .A1(_00203_),
    .S(mem_la_wdata[3]),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _25171_ (.A0(_00204_),
    .A1(_00220_),
    .S(mem_la_wdata[4]),
    .X(_13010_));
 sky130_fd_sc_hd__mux2_1 _25172_ (.A0(_00161_),
    .A1(_00163_),
    .S(mem_la_wdata[1]),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _25173_ (.A0(_00221_),
    .A1(_00222_),
    .S(mem_la_wdata[2]),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _25174_ (.A0(_00223_),
    .A1(_00226_),
    .S(mem_la_wdata[3]),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _25175_ (.A0(_00227_),
    .A1(_00234_),
    .S(mem_la_wdata[4]),
    .X(_13021_));
 sky130_fd_sc_hd__mux2_1 _25176_ (.A0(_00191_),
    .A1(_00193_),
    .S(mem_la_wdata[1]),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _25177_ (.A0(_00235_),
    .A1(_00236_),
    .S(mem_la_wdata[2]),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _25178_ (.A0(_00237_),
    .A1(_00240_),
    .S(mem_la_wdata[3]),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _25179_ (.A0(_00241_),
    .A1(_00248_),
    .S(mem_la_wdata[4]),
    .X(_13024_));
 sky130_fd_sc_hd__mux2_1 _25180_ (.A0(_00165_),
    .A1(_00169_),
    .S(mem_la_wdata[2]),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _25181_ (.A0(_00249_),
    .A1(_00250_),
    .S(mem_la_wdata[3]),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _25182_ (.A0(_00251_),
    .A1(_00254_),
    .S(mem_la_wdata[4]),
    .X(_13025_));
 sky130_fd_sc_hd__mux2_1 _25183_ (.A0(_00195_),
    .A1(_00199_),
    .S(mem_la_wdata[2]),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _25184_ (.A0(_00255_),
    .A1(_00256_),
    .S(mem_la_wdata[3]),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _25185_ (.A0(_00257_),
    .A1(_00260_),
    .S(mem_la_wdata[4]),
    .X(_13026_));
 sky130_fd_sc_hd__mux2_1 _25186_ (.A0(_00222_),
    .A1(_00224_),
    .S(mem_la_wdata[2]),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _25187_ (.A0(_00261_),
    .A1(_00262_),
    .S(mem_la_wdata[3]),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _25188_ (.A0(_00263_),
    .A1(_00266_),
    .S(mem_la_wdata[4]),
    .X(_13027_));
 sky130_fd_sc_hd__mux2_1 _25189_ (.A0(_00236_),
    .A1(_00238_),
    .S(mem_la_wdata[2]),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _25190_ (.A0(_00267_),
    .A1(_00268_),
    .S(mem_la_wdata[3]),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _25191_ (.A0(_00269_),
    .A1(_00272_),
    .S(mem_la_wdata[4]),
    .X(_13028_));
 sky130_fd_sc_hd__mux2_1 _25192_ (.A0(_00173_),
    .A1(_00181_),
    .S(mem_la_wdata[3]),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _25193_ (.A0(_00273_),
    .A1(_00274_),
    .S(mem_la_wdata[4]),
    .X(_13029_));
 sky130_fd_sc_hd__mux2_1 _25194_ (.A0(_00203_),
    .A1(_00211_),
    .S(mem_la_wdata[3]),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _25195_ (.A0(_00275_),
    .A1(_00276_),
    .S(mem_la_wdata[4]),
    .X(_13030_));
 sky130_fd_sc_hd__mux2_1 _25196_ (.A0(_00226_),
    .A1(_00230_),
    .S(mem_la_wdata[3]),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _25197_ (.A0(_00277_),
    .A1(_00278_),
    .S(mem_la_wdata[4]),
    .X(_13000_));
 sky130_fd_sc_hd__mux2_1 _25198_ (.A0(_00240_),
    .A1(_00244_),
    .S(mem_la_wdata[3]),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _25199_ (.A0(_00279_),
    .A1(_00280_),
    .S(mem_la_wdata[4]),
    .X(_13001_));
 sky130_fd_sc_hd__mux2_1 _25200_ (.A0(_00250_),
    .A1(_00252_),
    .S(mem_la_wdata[3]),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _25201_ (.A0(_00281_),
    .A1(_00282_),
    .S(mem_la_wdata[4]),
    .X(_13002_));
 sky130_fd_sc_hd__mux2_1 _25202_ (.A0(_00256_),
    .A1(_00258_),
    .S(mem_la_wdata[3]),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _25203_ (.A0(_00283_),
    .A1(_00284_),
    .S(mem_la_wdata[4]),
    .X(_13003_));
 sky130_fd_sc_hd__mux2_1 _25204_ (.A0(_00262_),
    .A1(_00264_),
    .S(mem_la_wdata[3]),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _25205_ (.A0(_00285_),
    .A1(_00286_),
    .S(mem_la_wdata[4]),
    .X(_13004_));
 sky130_fd_sc_hd__mux2_1 _25206_ (.A0(_00268_),
    .A1(_00270_),
    .S(mem_la_wdata[3]),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _25207_ (.A0(_00287_),
    .A1(_00288_),
    .S(mem_la_wdata[4]),
    .X(_13005_));
 sky130_fd_sc_hd__mux2_1 _25208_ (.A0(_00189_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13006_));
 sky130_fd_sc_hd__mux2_1 _25209_ (.A0(_00220_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13007_));
 sky130_fd_sc_hd__mux2_1 _25210_ (.A0(_00234_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13008_));
 sky130_fd_sc_hd__mux2_1 _25211_ (.A0(_00248_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13009_));
 sky130_fd_sc_hd__mux2_1 _25212_ (.A0(_00254_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13011_));
 sky130_fd_sc_hd__mux2_1 _25213_ (.A0(_00260_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13012_));
 sky130_fd_sc_hd__mux2_1 _25214_ (.A0(_00266_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13013_));
 sky130_fd_sc_hd__mux2_1 _25215_ (.A0(_00272_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13014_));
 sky130_fd_sc_hd__mux2_1 _25216_ (.A0(_00274_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13015_));
 sky130_fd_sc_hd__mux2_1 _25217_ (.A0(_00276_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13016_));
 sky130_fd_sc_hd__mux2_1 _25218_ (.A0(_00278_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13017_));
 sky130_fd_sc_hd__mux2_1 _25219_ (.A0(_00280_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13018_));
 sky130_fd_sc_hd__mux2_1 _25220_ (.A0(_00282_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13019_));
 sky130_fd_sc_hd__mux2_1 _25221_ (.A0(_00284_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13020_));
 sky130_fd_sc_hd__mux2_1 _25222_ (.A0(_00286_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13022_));
 sky130_fd_sc_hd__mux2_1 _25223_ (.A0(_00288_),
    .A1(_00216_),
    .S(mem_la_wdata[4]),
    .X(_13023_));
 sky130_fd_sc_hd__mux2_1 _25224_ (.A0(_01697_),
    .A1(_01698_),
    .S(\irq_state[1] ),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _25225_ (.A0(_01705_),
    .A1(_01699_),
    .S(_01700_),
    .X(_12982_));
 sky130_fd_sc_hd__mux2_1 _25226_ (.A0(_01720_),
    .A1(\irq_pending[0] ),
    .S(_01706_),
    .X(_12948_));
 sky130_fd_sc_hd__mux2_1 _25227_ (.A0(_01733_),
    .A1(\irq_pending[1] ),
    .S(_01706_),
    .X(_12959_));
 sky130_fd_sc_hd__mux2_1 _25228_ (.A0(_01746_),
    .A1(\irq_pending[2] ),
    .S(_01706_),
    .X(_12970_));
 sky130_fd_sc_hd__mux2_1 _25229_ (.A0(_01759_),
    .A1(\irq_pending[3] ),
    .S(_01706_),
    .X(_12973_));
 sky130_fd_sc_hd__mux2_1 _25230_ (.A0(_01772_),
    .A1(\irq_pending[4] ),
    .S(_01706_),
    .X(_12974_));
 sky130_fd_sc_hd__mux2_1 _25231_ (.A0(_01785_),
    .A1(\irq_pending[5] ),
    .S(_01706_),
    .X(_12975_));
 sky130_fd_sc_hd__mux2_1 _25232_ (.A0(_01798_),
    .A1(\irq_pending[6] ),
    .S(_01706_),
    .X(_12976_));
 sky130_fd_sc_hd__mux2_1 _25233_ (.A0(_01811_),
    .A1(\irq_pending[7] ),
    .S(_01706_),
    .X(_12977_));
 sky130_fd_sc_hd__mux2_1 _25234_ (.A0(_01825_),
    .A1(\irq_pending[8] ),
    .S(_01706_),
    .X(_12978_));
 sky130_fd_sc_hd__mux2_1 _25235_ (.A0(_01838_),
    .A1(\irq_pending[9] ),
    .S(_01706_),
    .X(_12979_));
 sky130_fd_sc_hd__mux2_1 _25236_ (.A0(_01851_),
    .A1(\irq_pending[10] ),
    .S(_01706_),
    .X(_12949_));
 sky130_fd_sc_hd__mux2_1 _25237_ (.A0(_01864_),
    .A1(\irq_pending[11] ),
    .S(_01706_),
    .X(_12950_));
 sky130_fd_sc_hd__mux2_1 _25238_ (.A0(_01877_),
    .A1(\irq_pending[12] ),
    .S(_01706_),
    .X(_12951_));
 sky130_fd_sc_hd__mux2_1 _25239_ (.A0(_01890_),
    .A1(\irq_pending[13] ),
    .S(_01706_),
    .X(_12952_));
 sky130_fd_sc_hd__mux2_1 _25240_ (.A0(_01903_),
    .A1(\irq_pending[14] ),
    .S(_01706_),
    .X(_12953_));
 sky130_fd_sc_hd__mux2_1 _25241_ (.A0(_01916_),
    .A1(\irq_pending[15] ),
    .S(_01706_),
    .X(_12954_));
 sky130_fd_sc_hd__mux2_1 _25242_ (.A0(_01925_),
    .A1(\irq_pending[16] ),
    .S(_01706_),
    .X(_12955_));
 sky130_fd_sc_hd__mux2_1 _25243_ (.A0(_01934_),
    .A1(\irq_pending[17] ),
    .S(_01706_),
    .X(_12956_));
 sky130_fd_sc_hd__mux2_1 _25244_ (.A0(_01943_),
    .A1(\irq_pending[18] ),
    .S(_01706_),
    .X(_12957_));
 sky130_fd_sc_hd__mux2_1 _25245_ (.A0(_01952_),
    .A1(\irq_pending[19] ),
    .S(_01706_),
    .X(_12958_));
 sky130_fd_sc_hd__mux2_1 _25246_ (.A0(_01961_),
    .A1(\irq_pending[20] ),
    .S(_01706_),
    .X(_12960_));
 sky130_fd_sc_hd__mux2_1 _25247_ (.A0(_01970_),
    .A1(\irq_pending[21] ),
    .S(_01706_),
    .X(_12961_));
 sky130_fd_sc_hd__mux2_1 _25248_ (.A0(_01979_),
    .A1(\irq_pending[22] ),
    .S(_01706_),
    .X(_12962_));
 sky130_fd_sc_hd__mux2_1 _25249_ (.A0(_01988_),
    .A1(\irq_pending[23] ),
    .S(_01706_),
    .X(_12963_));
 sky130_fd_sc_hd__mux2_1 _25250_ (.A0(_01997_),
    .A1(\irq_pending[24] ),
    .S(_01706_),
    .X(_12964_));
 sky130_fd_sc_hd__mux2_1 _25251_ (.A0(_02006_),
    .A1(\irq_pending[25] ),
    .S(_01706_),
    .X(_12965_));
 sky130_fd_sc_hd__mux2_1 _25252_ (.A0(_02015_),
    .A1(\irq_pending[26] ),
    .S(_01706_),
    .X(_12966_));
 sky130_fd_sc_hd__mux2_1 _25253_ (.A0(_02024_),
    .A1(\irq_pending[27] ),
    .S(_01706_),
    .X(_12967_));
 sky130_fd_sc_hd__mux2_1 _25254_ (.A0(_02033_),
    .A1(\irq_pending[28] ),
    .S(_01706_),
    .X(_12968_));
 sky130_fd_sc_hd__mux2_1 _25255_ (.A0(_02042_),
    .A1(\irq_pending[29] ),
    .S(_01706_),
    .X(_12969_));
 sky130_fd_sc_hd__mux2_1 _25256_ (.A0(_02051_),
    .A1(\irq_pending[30] ),
    .S(_01706_),
    .X(_12971_));
 sky130_fd_sc_hd__mux2_1 _25257_ (.A0(_02060_),
    .A1(\irq_pending[31] ),
    .S(_01706_),
    .X(_12972_));
 sky130_fd_sc_hd__mux2_1 _25258_ (.A0(_02061_),
    .A1(\cpu_state[2] ),
    .S(_02542_),
    .X(_12943_));
 sky130_fd_sc_hd__mux2_1 _25259_ (.A0(\decoded_rd[0] ),
    .A1(\irq_state[0] ),
    .S(_00308_),
    .X(_12942_));
 sky130_fd_sc_hd__mux2_1 _25260_ (.A0(_02062_),
    .A1(_02065_),
    .S(_02542_),
    .X(_12980_));
 sky130_fd_sc_hd__mux2_1 _25261_ (.A0(_02068_),
    .A1(_02066_),
    .S(_02067_),
    .X(_12981_));
 sky130_fd_sc_hd__mux2_1 _25262_ (.A0(_02166_),
    .A1(_00291_),
    .S(_00290_),
    .X(_12944_));
 sky130_fd_sc_hd__mux2_1 _25263_ (.A0(_02166_),
    .A1(mem_do_wdata),
    .S(_00290_),
    .X(_12945_));
 sky130_fd_sc_hd__mux2_1 _25264_ (.A0(_00271_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _25265_ (.A0(_00265_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _25266_ (.A0(_00259_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _25267_ (.A0(_00253_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _25268_ (.A0(_00247_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _25269_ (.A0(_00233_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _25270_ (.A0(_00219_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _25271_ (.A0(_00188_),
    .A1(_00216_),
    .S(mem_la_wdata[3]),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _25272_ (.A0(_00270_),
    .A1(_00271_),
    .S(mem_la_wdata[3]),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _25273_ (.A0(_00246_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _25274_ (.A0(_00243_),
    .A1(_00245_),
    .S(mem_la_wdata[2]),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _25275_ (.A0(_00239_),
    .A1(_00242_),
    .S(mem_la_wdata[2]),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _25276_ (.A0(_00264_),
    .A1(_00265_),
    .S(mem_la_wdata[3]),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _25277_ (.A0(_00232_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _25278_ (.A0(_00229_),
    .A1(_00231_),
    .S(mem_la_wdata[2]),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _25279_ (.A0(_00225_),
    .A1(_00228_),
    .S(mem_la_wdata[2]),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _25280_ (.A0(_00258_),
    .A1(_00259_),
    .S(mem_la_wdata[3]),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _25281_ (.A0(_00218_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _25282_ (.A0(_00210_),
    .A1(_00214_),
    .S(mem_la_wdata[2]),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _25283_ (.A0(_00202_),
    .A1(_00207_),
    .S(mem_la_wdata[2]),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _25284_ (.A0(_00252_),
    .A1(_00253_),
    .S(mem_la_wdata[3]),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _25285_ (.A0(_00187_),
    .A1(_00216_),
    .S(mem_la_wdata[2]),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _25286_ (.A0(_00180_),
    .A1(_00184_),
    .S(mem_la_wdata[2]),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _25287_ (.A0(_00172_),
    .A1(_00177_),
    .S(mem_la_wdata[2]),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _25288_ (.A0(_00244_),
    .A1(_00247_),
    .S(mem_la_wdata[3]),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _25289_ (.A0(_00245_),
    .A1(_00246_),
    .S(mem_la_wdata[2]),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _25290_ (.A0(_00217_),
    .A1(_00216_),
    .S(mem_la_wdata[1]),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _25291_ (.A0(_00213_),
    .A1(_00215_),
    .S(mem_la_wdata[1]),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _25292_ (.A0(_00242_),
    .A1(_00243_),
    .S(mem_la_wdata[2]),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _25293_ (.A0(_00209_),
    .A1(_00212_),
    .S(mem_la_wdata[1]),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _25294_ (.A0(_00206_),
    .A1(_00208_),
    .S(mem_la_wdata[1]),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _25295_ (.A0(_00238_),
    .A1(_00239_),
    .S(mem_la_wdata[2]),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _25296_ (.A0(_00201_),
    .A1(_00205_),
    .S(mem_la_wdata[1]),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _25297_ (.A0(_00198_),
    .A1(_00200_),
    .S(mem_la_wdata[1]),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _25298_ (.A0(_00194_),
    .A1(_00197_),
    .S(mem_la_wdata[1]),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _25299_ (.A0(_00230_),
    .A1(_00233_),
    .S(mem_la_wdata[3]),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _25300_ (.A0(_00231_),
    .A1(_00232_),
    .S(mem_la_wdata[2]),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _25301_ (.A0(_00186_),
    .A1(_00216_),
    .S(mem_la_wdata[1]),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _25302_ (.A0(_00183_),
    .A1(_00185_),
    .S(mem_la_wdata[1]),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _25303_ (.A0(_00228_),
    .A1(_00229_),
    .S(mem_la_wdata[2]),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _25304_ (.A0(_00179_),
    .A1(_00182_),
    .S(mem_la_wdata[1]),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _25305_ (.A0(_00176_),
    .A1(_00178_),
    .S(mem_la_wdata[1]),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _25306_ (.A0(_00224_),
    .A1(_00225_),
    .S(mem_la_wdata[2]),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _25307_ (.A0(_00171_),
    .A1(_00175_),
    .S(mem_la_wdata[1]),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _25308_ (.A0(_00168_),
    .A1(_00170_),
    .S(mem_la_wdata[1]),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _25309_ (.A0(_00164_),
    .A1(_00167_),
    .S(mem_la_wdata[1]),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _25310_ (.A0(_00211_),
    .A1(_00219_),
    .S(mem_la_wdata[3]),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _25311_ (.A0(_00214_),
    .A1(_00218_),
    .S(mem_la_wdata[2]),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _25312_ (.A0(_00215_),
    .A1(_00217_),
    .S(mem_la_wdata[1]),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _25313_ (.A0(pcpi_rs1[31]),
    .A1(_00216_),
    .S(mem_la_wdata[0]),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _25314_ (.A0(pcpi_rs1[29]),
    .A1(pcpi_rs1[30]),
    .S(mem_la_wdata[0]),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _25315_ (.A0(_00212_),
    .A1(_00213_),
    .S(mem_la_wdata[1]),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _25316_ (.A0(pcpi_rs1[27]),
    .A1(pcpi_rs1[28]),
    .S(mem_la_wdata[0]),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _25317_ (.A0(pcpi_rs1[25]),
    .A1(pcpi_rs1[26]),
    .S(mem_la_wdata[0]),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _25318_ (.A0(_00207_),
    .A1(_00210_),
    .S(mem_la_wdata[2]),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _25319_ (.A0(_00208_),
    .A1(_00209_),
    .S(mem_la_wdata[1]),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _25320_ (.A0(pcpi_rs1[23]),
    .A1(pcpi_rs1[24]),
    .S(mem_la_wdata[0]),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _25321_ (.A0(pcpi_rs1[21]),
    .A1(pcpi_rs1[22]),
    .S(mem_la_wdata[0]),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _25322_ (.A0(_00205_),
    .A1(_00206_),
    .S(mem_la_wdata[1]),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _25323_ (.A0(pcpi_rs1[19]),
    .A1(pcpi_rs1[20]),
    .S(mem_la_wdata[0]),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _25324_ (.A0(pcpi_rs1[17]),
    .A1(pcpi_rs1[18]),
    .S(mem_la_wdata[0]),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _25325_ (.A0(_00199_),
    .A1(_00202_),
    .S(mem_la_wdata[2]),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _25326_ (.A0(_00200_),
    .A1(_00201_),
    .S(mem_la_wdata[1]),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _25327_ (.A0(pcpi_rs1[15]),
    .A1(pcpi_rs1[16]),
    .S(mem_la_wdata[0]),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _25328_ (.A0(pcpi_rs1[13]),
    .A1(pcpi_rs1[14]),
    .S(mem_la_wdata[0]),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _25329_ (.A0(_00197_),
    .A1(_00198_),
    .S(mem_la_wdata[1]),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _25330_ (.A0(pcpi_rs1[11]),
    .A1(pcpi_rs1[12]),
    .S(mem_la_wdata[0]),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _25331_ (.A0(pcpi_rs1[9]),
    .A1(pcpi_rs1[10]),
    .S(mem_la_wdata[0]),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _25332_ (.A0(_00193_),
    .A1(_00194_),
    .S(mem_la_wdata[1]),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _25333_ (.A0(pcpi_rs1[7]),
    .A1(pcpi_rs1[8]),
    .S(mem_la_wdata[0]),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _25334_ (.A0(pcpi_rs1[5]),
    .A1(pcpi_rs1[6]),
    .S(mem_la_wdata[0]),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _25335_ (.A0(pcpi_rs1[3]),
    .A1(pcpi_rs1[4]),
    .S(mem_la_wdata[0]),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _25336_ (.A0(_00181_),
    .A1(_00188_),
    .S(mem_la_wdata[3]),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _25337_ (.A0(_00184_),
    .A1(_00187_),
    .S(mem_la_wdata[2]),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _25338_ (.A0(_00185_),
    .A1(_00186_),
    .S(mem_la_wdata[1]),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _25339_ (.A0(pcpi_rs1[30]),
    .A1(pcpi_rs1[31]),
    .S(mem_la_wdata[0]),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _25340_ (.A0(pcpi_rs1[28]),
    .A1(pcpi_rs1[29]),
    .S(mem_la_wdata[0]),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _25341_ (.A0(_00182_),
    .A1(_00183_),
    .S(mem_la_wdata[1]),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _25342_ (.A0(pcpi_rs1[26]),
    .A1(pcpi_rs1[27]),
    .S(mem_la_wdata[0]),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _25343_ (.A0(pcpi_rs1[24]),
    .A1(pcpi_rs1[25]),
    .S(mem_la_wdata[0]),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _25344_ (.A0(_00177_),
    .A1(_00180_),
    .S(mem_la_wdata[2]),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _25345_ (.A0(_00178_),
    .A1(_00179_),
    .S(mem_la_wdata[1]),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _25346_ (.A0(pcpi_rs1[22]),
    .A1(pcpi_rs1[23]),
    .S(mem_la_wdata[0]),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _25347_ (.A0(pcpi_rs1[20]),
    .A1(pcpi_rs1[21]),
    .S(mem_la_wdata[0]),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _25348_ (.A0(_00175_),
    .A1(_00176_),
    .S(mem_la_wdata[1]),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _25349_ (.A0(pcpi_rs1[18]),
    .A1(pcpi_rs1[19]),
    .S(mem_la_wdata[0]),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _25350_ (.A0(pcpi_rs1[16]),
    .A1(pcpi_rs1[17]),
    .S(mem_la_wdata[0]),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _25351_ (.A0(_00169_),
    .A1(_00172_),
    .S(mem_la_wdata[2]),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _25352_ (.A0(_00170_),
    .A1(_00171_),
    .S(mem_la_wdata[1]),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _25353_ (.A0(pcpi_rs1[14]),
    .A1(pcpi_rs1[15]),
    .S(mem_la_wdata[0]),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _25354_ (.A0(pcpi_rs1[12]),
    .A1(pcpi_rs1[13]),
    .S(mem_la_wdata[0]),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _25355_ (.A0(_00167_),
    .A1(_00168_),
    .S(mem_la_wdata[1]),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _25356_ (.A0(pcpi_rs1[10]),
    .A1(pcpi_rs1[11]),
    .S(mem_la_wdata[0]),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _25357_ (.A0(pcpi_rs1[8]),
    .A1(pcpi_rs1[9]),
    .S(mem_la_wdata[0]),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _25358_ (.A0(_00163_),
    .A1(_00164_),
    .S(mem_la_wdata[1]),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _25359_ (.A0(pcpi_rs1[6]),
    .A1(pcpi_rs1[7]),
    .S(mem_la_wdata[0]),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _25360_ (.A0(pcpi_rs1[4]),
    .A1(pcpi_rs1[5]),
    .S(mem_la_wdata[0]),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _25361_ (.A0(pcpi_rs1[2]),
    .A1(pcpi_rs1[3]),
    .S(mem_la_wdata[0]),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _25362_ (.A0(pcpi_rs1[29]),
    .A1(pcpi_rs1[28]),
    .S(mem_la_wdata[0]),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _25363_ (.A0(pcpi_rs1[28]),
    .A1(pcpi_rs1[27]),
    .S(mem_la_wdata[0]),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _25364_ (.A0(_00140_),
    .A1(_00132_),
    .S(mem_la_wdata[1]),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _25365_ (.A0(pcpi_rs1[27]),
    .A1(pcpi_rs1[26]),
    .S(mem_la_wdata[0]),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _25366_ (.A0(_00136_),
    .A1(_00128_),
    .S(mem_la_wdata[1]),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _25367_ (.A0(pcpi_rs1[26]),
    .A1(pcpi_rs1[25]),
    .S(mem_la_wdata[0]),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _25368_ (.A0(_00132_),
    .A1(_00123_),
    .S(mem_la_wdata[1]),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _25369_ (.A0(pcpi_rs1[25]),
    .A1(pcpi_rs1[24]),
    .S(mem_la_wdata[0]),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _25370_ (.A0(_00128_),
    .A1(_00117_),
    .S(mem_la_wdata[1]),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _25371_ (.A0(pcpi_rs1[24]),
    .A1(pcpi_rs1[23]),
    .S(mem_la_wdata[0]),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _25372_ (.A0(_00098_),
    .A1(_00100_),
    .S(mem_la_wdata[2]),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _25373_ (.A0(_00124_),
    .A1(_00097_),
    .S(mem_la_wdata[2]),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _25374_ (.A0(_00123_),
    .A1(_00111_),
    .S(mem_la_wdata[1]),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _25375_ (.A0(pcpi_rs1[23]),
    .A1(pcpi_rs1[22]),
    .S(mem_la_wdata[0]),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _25376_ (.A0(_00101_),
    .A1(_00094_),
    .S(mem_la_wdata[2]),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _25377_ (.A0(_00088_),
    .A1(_00090_),
    .S(mem_la_wdata[2]),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _25378_ (.A0(_00118_),
    .A1(_00087_),
    .S(mem_la_wdata[2]),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _25379_ (.A0(_00117_),
    .A1(_00105_),
    .S(mem_la_wdata[1]),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _25380_ (.A0(pcpi_rs1[22]),
    .A1(pcpi_rs1[21]),
    .S(mem_la_wdata[0]),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _25381_ (.A0(_00091_),
    .A1(_00084_),
    .S(mem_la_wdata[2]),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _25382_ (.A0(_00074_),
    .A1(_00078_),
    .S(mem_la_wdata[2]),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _25383_ (.A0(_00112_),
    .A1(_00071_),
    .S(mem_la_wdata[2]),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _25384_ (.A0(_00111_),
    .A1(_00096_),
    .S(mem_la_wdata[1]),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _25385_ (.A0(pcpi_rs1[21]),
    .A1(pcpi_rs1[20]),
    .S(mem_la_wdata[0]),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _25386_ (.A0(_00081_),
    .A1(_00067_),
    .S(mem_la_wdata[2]),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _25387_ (.A0(_00056_),
    .A1(_00060_),
    .S(mem_la_wdata[2]),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _25388_ (.A0(_00106_),
    .A1(_00053_),
    .S(mem_la_wdata[2]),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _25389_ (.A0(_00105_),
    .A1(_00086_),
    .S(mem_la_wdata[1]),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _25390_ (.A0(pcpi_rs1[20]),
    .A1(pcpi_rs1[19]),
    .S(mem_la_wdata[0]),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _25391_ (.A0(_00063_),
    .A1(_00049_),
    .S(mem_la_wdata[2]),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _25392_ (.A0(_00100_),
    .A1(_00101_),
    .S(mem_la_wdata[2]),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _25393_ (.A0(_00077_),
    .A1(_00079_),
    .S(mem_la_wdata[1]),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _25394_ (.A0(_00073_),
    .A1(_00076_),
    .S(mem_la_wdata[1]),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _25395_ (.A0(_00097_),
    .A1(_00098_),
    .S(mem_la_wdata[2]),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _25396_ (.A0(_00070_),
    .A1(_00072_),
    .S(mem_la_wdata[1]),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _25397_ (.A0(_00096_),
    .A1(_00069_),
    .S(mem_la_wdata[1]),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _25398_ (.A0(pcpi_rs1[19]),
    .A1(pcpi_rs1[18]),
    .S(mem_la_wdata[0]),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _25399_ (.A0(_00080_),
    .A1(_00066_),
    .S(mem_la_wdata[1]),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _25400_ (.A0(_00090_),
    .A1(_00091_),
    .S(mem_la_wdata[2]),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _25401_ (.A0(_00059_),
    .A1(_00061_),
    .S(mem_la_wdata[1]),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _25402_ (.A0(_00055_),
    .A1(_00058_),
    .S(mem_la_wdata[1]),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _25403_ (.A0(_00087_),
    .A1(_00088_),
    .S(mem_la_wdata[2]),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _25404_ (.A0(_00052_),
    .A1(_00054_),
    .S(mem_la_wdata[1]),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _25405_ (.A0(_00086_),
    .A1(_00051_),
    .S(mem_la_wdata[1]),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _25406_ (.A0(pcpi_rs1[18]),
    .A1(pcpi_rs1[17]),
    .S(mem_la_wdata[0]),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _25407_ (.A0(_00062_),
    .A1(_00048_),
    .S(mem_la_wdata[1]),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _25408_ (.A0(_00078_),
    .A1(_00081_),
    .S(mem_la_wdata[2]),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _25409_ (.A0(_00079_),
    .A1(_00080_),
    .S(mem_la_wdata[1]),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _25410_ (.A0(pcpi_rs1[3]),
    .A1(pcpi_rs1[2]),
    .S(mem_la_wdata[0]),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _25411_ (.A0(pcpi_rs1[5]),
    .A1(pcpi_rs1[4]),
    .S(mem_la_wdata[0]),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _25412_ (.A0(_00076_),
    .A1(_00077_),
    .S(mem_la_wdata[1]),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _25413_ (.A0(pcpi_rs1[7]),
    .A1(pcpi_rs1[6]),
    .S(mem_la_wdata[0]),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _25414_ (.A0(pcpi_rs1[9]),
    .A1(pcpi_rs1[8]),
    .S(mem_la_wdata[0]),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _25415_ (.A0(_00071_),
    .A1(_00074_),
    .S(mem_la_wdata[2]),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _25416_ (.A0(_00072_),
    .A1(_00073_),
    .S(mem_la_wdata[1]),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _25417_ (.A0(pcpi_rs1[11]),
    .A1(pcpi_rs1[10]),
    .S(mem_la_wdata[0]),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _25418_ (.A0(pcpi_rs1[13]),
    .A1(pcpi_rs1[12]),
    .S(mem_la_wdata[0]),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _25419_ (.A0(_00069_),
    .A1(_00070_),
    .S(mem_la_wdata[1]),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _25420_ (.A0(pcpi_rs1[15]),
    .A1(pcpi_rs1[14]),
    .S(mem_la_wdata[0]),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _25421_ (.A0(pcpi_rs1[17]),
    .A1(pcpi_rs1[16]),
    .S(mem_la_wdata[0]),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _25422_ (.A0(pcpi_rs1[1]),
    .A1(pcpi_rs1[0]),
    .S(mem_la_wdata[0]),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _25423_ (.A0(_00060_),
    .A1(_00063_),
    .S(mem_la_wdata[2]),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _25424_ (.A0(_00061_),
    .A1(_00062_),
    .S(mem_la_wdata[1]),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _25425_ (.A0(pcpi_rs1[2]),
    .A1(pcpi_rs1[1]),
    .S(mem_la_wdata[0]),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _25426_ (.A0(pcpi_rs1[4]),
    .A1(pcpi_rs1[3]),
    .S(mem_la_wdata[0]),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _25427_ (.A0(_00058_),
    .A1(_00059_),
    .S(mem_la_wdata[1]),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _25428_ (.A0(pcpi_rs1[6]),
    .A1(pcpi_rs1[5]),
    .S(mem_la_wdata[0]),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _25429_ (.A0(pcpi_rs1[8]),
    .A1(pcpi_rs1[7]),
    .S(mem_la_wdata[0]),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _25430_ (.A0(_00053_),
    .A1(_00056_),
    .S(mem_la_wdata[2]),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _25431_ (.A0(_00054_),
    .A1(_00055_),
    .S(mem_la_wdata[1]),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _25432_ (.A0(pcpi_rs1[10]),
    .A1(pcpi_rs1[9]),
    .S(mem_la_wdata[0]),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _25433_ (.A0(pcpi_rs1[12]),
    .A1(pcpi_rs1[11]),
    .S(mem_la_wdata[0]),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _25434_ (.A0(_00051_),
    .A1(_00052_),
    .S(mem_la_wdata[1]),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _25435_ (.A0(pcpi_rs1[14]),
    .A1(pcpi_rs1[13]),
    .S(mem_la_wdata[0]),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _25436_ (.A0(pcpi_rs1[16]),
    .A1(pcpi_rs1[15]),
    .S(mem_la_wdata[0]),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _25437_ (.A0(_02408_),
    .A1(pcpi_rs2[31]),
    .S(instr_sub),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _25438_ (.A0(_02406_),
    .A1(_02405_),
    .S(instr_sub),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _25439_ (.A0(_02403_),
    .A1(_02402_),
    .S(instr_sub),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _25440_ (.A0(_02400_),
    .A1(_02399_),
    .S(instr_sub),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _25441_ (.A0(_02397_),
    .A1(_02396_),
    .S(instr_sub),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _25442_ (.A0(_02394_),
    .A1(_02393_),
    .S(instr_sub),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _25443_ (.A0(_02391_),
    .A1(_02390_),
    .S(instr_sub),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _25444_ (.A0(_02388_),
    .A1(_02387_),
    .S(instr_sub),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _25445_ (.A0(_02385_),
    .A1(_02384_),
    .S(instr_sub),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _25446_ (.A0(_02382_),
    .A1(_02381_),
    .S(instr_sub),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _25447_ (.A0(_02379_),
    .A1(_02378_),
    .S(instr_sub),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _25448_ (.A0(_02376_),
    .A1(_02375_),
    .S(instr_sub),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _25449_ (.A0(_02373_),
    .A1(_02372_),
    .S(instr_sub),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_1 _25450_ (.A0(_02370_),
    .A1(_02369_),
    .S(instr_sub),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _25451_ (.A0(_02367_),
    .A1(_02366_),
    .S(instr_sub),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_1 _25452_ (.A0(_02364_),
    .A1(_02363_),
    .S(instr_sub),
    .X(_02365_));
 sky130_fd_sc_hd__mux2_1 _25453_ (.A0(_02361_),
    .A1(_02360_),
    .S(instr_sub),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _25454_ (.A0(_02358_),
    .A1(_02357_),
    .S(instr_sub),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _25455_ (.A0(_02355_),
    .A1(_02354_),
    .S(instr_sub),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _25456_ (.A0(_02352_),
    .A1(_02351_),
    .S(instr_sub),
    .X(_02353_));
 sky130_fd_sc_hd__mux2_1 _25457_ (.A0(_02349_),
    .A1(_02348_),
    .S(instr_sub),
    .X(_02350_));
 sky130_fd_sc_hd__mux2_1 _25458_ (.A0(_02346_),
    .A1(_02345_),
    .S(instr_sub),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_1 _25459_ (.A0(_02343_),
    .A1(_02342_),
    .S(instr_sub),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_1 _25460_ (.A0(_02340_),
    .A1(_02339_),
    .S(instr_sub),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _25461_ (.A0(_02337_),
    .A1(_02336_),
    .S(instr_sub),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _25462_ (.A0(_02334_),
    .A1(_02333_),
    .S(instr_sub),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _25463_ (.A0(_02331_),
    .A1(_02330_),
    .S(instr_sub),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _25464_ (.A0(_02328_),
    .A1(_02327_),
    .S(instr_sub),
    .X(_02329_));
 sky130_fd_sc_hd__mux2_1 _25465_ (.A0(_02325_),
    .A1(_02324_),
    .S(instr_sub),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _25466_ (.A0(_02322_),
    .A1(_02321_),
    .S(instr_sub),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _25467_ (.A0(_02319_),
    .A1(_02318_),
    .S(instr_sub),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _25468_ (.A0(_02313_),
    .A1(_02314_),
    .S(_00306_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _25469_ (.A0(_02311_),
    .A1(_02315_),
    .S(_00303_),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _25470_ (.A0(_02311_),
    .A1(_02312_),
    .S(_00305_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _25471_ (.A0(_02307_),
    .A1(_02308_),
    .S(\irq_state[1] ),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _25472_ (.A0(_02309_),
    .A1(_02307_),
    .S(_02217_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _25473_ (.A0(_02302_),
    .A1(\irq_pending[0] ),
    .S(_01208_),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _25474_ (.A0(\reg_out[0] ),
    .A1(\alu_out_q[0] ),
    .S(latched_stalu),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _25475_ (.A0(_02063_),
    .A1(_00343_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _25476_ (.A0(_02056_),
    .A1(_02055_),
    .S(_01714_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _25477_ (.A0(_02058_),
    .A1(_02057_),
    .S(_01717_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _25478_ (.A0(\pcpi_mul.rd[31] ),
    .A1(\pcpi_mul.rd[63] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _25479_ (.A0(_01908_),
    .A1(_02052_),
    .S(_01816_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _25480_ (.A0(_02047_),
    .A1(_02046_),
    .S(_01714_),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _25481_ (.A0(_02049_),
    .A1(_02048_),
    .S(_01717_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _25482_ (.A0(\pcpi_mul.rd[30] ),
    .A1(\pcpi_mul.rd[62] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _25483_ (.A0(_01908_),
    .A1(_02043_),
    .S(_01816_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _25484_ (.A0(_02038_),
    .A1(_02037_),
    .S(_01714_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _25485_ (.A0(_02040_),
    .A1(_02039_),
    .S(_01717_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _25486_ (.A0(\pcpi_mul.rd[29] ),
    .A1(\pcpi_mul.rd[61] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _25487_ (.A0(_01908_),
    .A1(_02034_),
    .S(_01816_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _25488_ (.A0(_02029_),
    .A1(_02028_),
    .S(_01714_),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_1 _25489_ (.A0(_02031_),
    .A1(_02030_),
    .S(_01717_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _25490_ (.A0(\pcpi_mul.rd[28] ),
    .A1(\pcpi_mul.rd[60] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_1 _25491_ (.A0(_01908_),
    .A1(_02025_),
    .S(_01816_),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _25492_ (.A0(_02020_),
    .A1(_02019_),
    .S(_01714_),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_1 _25493_ (.A0(_02022_),
    .A1(_02021_),
    .S(_01717_),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _25494_ (.A0(\pcpi_mul.rd[27] ),
    .A1(\pcpi_mul.rd[59] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _25495_ (.A0(_01908_),
    .A1(_02016_),
    .S(_01816_),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _25496_ (.A0(_02011_),
    .A1(_02010_),
    .S(_01714_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _25497_ (.A0(_02013_),
    .A1(_02012_),
    .S(_01717_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _25498_ (.A0(\pcpi_mul.rd[26] ),
    .A1(\pcpi_mul.rd[58] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _25499_ (.A0(_01908_),
    .A1(_02007_),
    .S(_01816_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _25500_ (.A0(_02002_),
    .A1(_02001_),
    .S(_01714_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_1 _25501_ (.A0(_02004_),
    .A1(_02003_),
    .S(_01717_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _25502_ (.A0(\pcpi_mul.rd[25] ),
    .A1(\pcpi_mul.rd[57] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_1 _25503_ (.A0(_01908_),
    .A1(_01998_),
    .S(_01816_),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _25504_ (.A0(_01993_),
    .A1(_01992_),
    .S(_01714_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_1 _25505_ (.A0(_01995_),
    .A1(_01994_),
    .S(_01717_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _25506_ (.A0(\pcpi_mul.rd[24] ),
    .A1(\pcpi_mul.rd[56] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _25507_ (.A0(_01908_),
    .A1(_01989_),
    .S(_01816_),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_1 _25508_ (.A0(_01984_),
    .A1(_01983_),
    .S(_01714_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _25509_ (.A0(_01986_),
    .A1(_01985_),
    .S(_01717_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _25510_ (.A0(\pcpi_mul.rd[23] ),
    .A1(\pcpi_mul.rd[55] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _25511_ (.A0(_01908_),
    .A1(_01980_),
    .S(_01816_),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _25512_ (.A0(_01975_),
    .A1(_01974_),
    .S(_01714_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_1 _25513_ (.A0(_01977_),
    .A1(_01976_),
    .S(_01717_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _25514_ (.A0(\pcpi_mul.rd[22] ),
    .A1(\pcpi_mul.rd[54] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _25515_ (.A0(_01908_),
    .A1(_01971_),
    .S(_01816_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _25516_ (.A0(_01966_),
    .A1(_01965_),
    .S(_01714_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _25517_ (.A0(_01968_),
    .A1(_01967_),
    .S(_01717_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _25518_ (.A0(\pcpi_mul.rd[21] ),
    .A1(\pcpi_mul.rd[53] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _25519_ (.A0(_01908_),
    .A1(_01962_),
    .S(_01816_),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _25520_ (.A0(_01957_),
    .A1(_01956_),
    .S(_01714_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_1 _25521_ (.A0(_01959_),
    .A1(_01958_),
    .S(_01717_),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_1 _25522_ (.A0(\pcpi_mul.rd[20] ),
    .A1(\pcpi_mul.rd[52] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _25523_ (.A0(_01908_),
    .A1(_01953_),
    .S(_01816_),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _25524_ (.A0(_01948_),
    .A1(_01947_),
    .S(_01714_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _25525_ (.A0(_01950_),
    .A1(_01949_),
    .S(_01717_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _25526_ (.A0(\pcpi_mul.rd[19] ),
    .A1(\pcpi_mul.rd[51] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _25527_ (.A0(_01908_),
    .A1(_01944_),
    .S(_01816_),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _25528_ (.A0(_01939_),
    .A1(_01938_),
    .S(_01714_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_1 _25529_ (.A0(_01941_),
    .A1(_01940_),
    .S(_01717_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _25530_ (.A0(\pcpi_mul.rd[18] ),
    .A1(\pcpi_mul.rd[50] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _25531_ (.A0(_01908_),
    .A1(_01935_),
    .S(_01816_),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_1 _25532_ (.A0(_01930_),
    .A1(_01929_),
    .S(_01714_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_1 _25533_ (.A0(_01932_),
    .A1(_01931_),
    .S(_01717_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _25534_ (.A0(\pcpi_mul.rd[17] ),
    .A1(\pcpi_mul.rd[49] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _25535_ (.A0(_01908_),
    .A1(_01926_),
    .S(_01816_),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _25536_ (.A0(_01921_),
    .A1(_01920_),
    .S(_01714_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_1 _25537_ (.A0(_01923_),
    .A1(_01922_),
    .S(_01717_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _25538_ (.A0(\pcpi_mul.rd[16] ),
    .A1(\pcpi_mul.rd[48] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _25539_ (.A0(_01908_),
    .A1(_01917_),
    .S(_01816_),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_1 _25540_ (.A0(_01912_),
    .A1(_01911_),
    .S(_01714_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _25541_ (.A0(_01914_),
    .A1(_01913_),
    .S(_01717_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _25542_ (.A0(\pcpi_mul.rd[15] ),
    .A1(\pcpi_mul.rd[47] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _25543_ (.A0(_01908_),
    .A1(_01907_),
    .S(_01816_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _25544_ (.A0(_01906_),
    .A1(_01904_),
    .S(_01683_),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _25545_ (.A0(mem_rdata[15]),
    .A1(mem_rdata[31]),
    .S(pcpi_rs1[1]),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _25546_ (.A0(_01899_),
    .A1(_01898_),
    .S(_01714_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_1 _25547_ (.A0(_01901_),
    .A1(_01900_),
    .S(_01717_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _25548_ (.A0(\pcpi_mul.rd[14] ),
    .A1(\pcpi_mul.rd[46] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _25549_ (.A0(_01895_),
    .A1(_01894_),
    .S(_01816_),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _25550_ (.A0(_01893_),
    .A1(_01891_),
    .S(_01683_),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _25551_ (.A0(mem_rdata[14]),
    .A1(mem_rdata[30]),
    .S(pcpi_rs1[1]),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _25552_ (.A0(_01886_),
    .A1(_01885_),
    .S(_01714_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _25553_ (.A0(_01888_),
    .A1(_01887_),
    .S(_01717_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _25554_ (.A0(\pcpi_mul.rd[13] ),
    .A1(\pcpi_mul.rd[45] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _25555_ (.A0(_01882_),
    .A1(_01881_),
    .S(_01816_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _25556_ (.A0(_01880_),
    .A1(_01878_),
    .S(_01683_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _25557_ (.A0(mem_rdata[13]),
    .A1(mem_rdata[29]),
    .S(pcpi_rs1[1]),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _25558_ (.A0(_01873_),
    .A1(_01872_),
    .S(_01714_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _25559_ (.A0(_01875_),
    .A1(_01874_),
    .S(_01717_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _25560_ (.A0(\pcpi_mul.rd[12] ),
    .A1(\pcpi_mul.rd[44] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _25561_ (.A0(_01869_),
    .A1(_01868_),
    .S(_01816_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _25562_ (.A0(_01867_),
    .A1(_01865_),
    .S(_01683_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _25563_ (.A0(mem_rdata[12]),
    .A1(mem_rdata[28]),
    .S(pcpi_rs1[1]),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _25564_ (.A0(_01860_),
    .A1(_01859_),
    .S(_01714_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _25565_ (.A0(_01862_),
    .A1(_01861_),
    .S(_01717_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _25566_ (.A0(\pcpi_mul.rd[11] ),
    .A1(\pcpi_mul.rd[43] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _25567_ (.A0(_01856_),
    .A1(_01855_),
    .S(_01816_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _25568_ (.A0(_01854_),
    .A1(_01852_),
    .S(_01683_),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _25569_ (.A0(mem_rdata[11]),
    .A1(mem_rdata[27]),
    .S(pcpi_rs1[1]),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _25570_ (.A0(_01847_),
    .A1(_01846_),
    .S(_01714_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _25571_ (.A0(_01849_),
    .A1(_01848_),
    .S(_01717_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _25572_ (.A0(\pcpi_mul.rd[10] ),
    .A1(\pcpi_mul.rd[42] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _25573_ (.A0(_01843_),
    .A1(_01842_),
    .S(_01816_),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _25574_ (.A0(_01841_),
    .A1(_01839_),
    .S(_01683_),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _25575_ (.A0(mem_rdata[10]),
    .A1(mem_rdata[26]),
    .S(pcpi_rs1[1]),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _25576_ (.A0(_01834_),
    .A1(_01833_),
    .S(_01714_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _25577_ (.A0(_01836_),
    .A1(_01835_),
    .S(_01717_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _25578_ (.A0(\pcpi_mul.rd[9] ),
    .A1(\pcpi_mul.rd[41] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _25579_ (.A0(_01830_),
    .A1(_01829_),
    .S(_01816_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _25580_ (.A0(_01828_),
    .A1(_01826_),
    .S(_01683_),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _25581_ (.A0(mem_rdata[9]),
    .A1(mem_rdata[25]),
    .S(pcpi_rs1[1]),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _25582_ (.A0(_01821_),
    .A1(_01820_),
    .S(_01714_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _25583_ (.A0(_01823_),
    .A1(_01822_),
    .S(_01717_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _25584_ (.A0(\pcpi_mul.rd[8] ),
    .A1(\pcpi_mul.rd[40] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _25585_ (.A0(_01817_),
    .A1(_01815_),
    .S(_01816_),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _25586_ (.A0(_01814_),
    .A1(_01812_),
    .S(_01683_),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _25587_ (.A0(mem_rdata[8]),
    .A1(mem_rdata[24]),
    .S(pcpi_rs1[1]),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _25588_ (.A0(_01807_),
    .A1(_01806_),
    .S(_01714_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _25589_ (.A0(_01809_),
    .A1(_01808_),
    .S(_01717_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _25590_ (.A0(\pcpi_mul.rd[7] ),
    .A1(\pcpi_mul.rd[39] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _25591_ (.A0(_01803_),
    .A1(_01799_),
    .S(_01683_),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _25592_ (.A0(mem_rdata[7]),
    .A1(mem_rdata[23]),
    .S(pcpi_rs1[1]),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _25593_ (.A0(_01800_),
    .A1(_01799_),
    .S(_00304_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _25594_ (.A0(_01794_),
    .A1(_01793_),
    .S(_01714_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _25595_ (.A0(_01796_),
    .A1(_01795_),
    .S(_01717_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _25596_ (.A0(\pcpi_mul.rd[6] ),
    .A1(\pcpi_mul.rd[38] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _25597_ (.A0(_01790_),
    .A1(_01786_),
    .S(_01683_),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _25598_ (.A0(mem_rdata[6]),
    .A1(mem_rdata[22]),
    .S(pcpi_rs1[1]),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _25599_ (.A0(_01787_),
    .A1(_01786_),
    .S(_00304_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _25600_ (.A0(_01781_),
    .A1(_01780_),
    .S(_01714_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _25601_ (.A0(_01783_),
    .A1(_01782_),
    .S(_01717_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _25602_ (.A0(\pcpi_mul.rd[5] ),
    .A1(\pcpi_mul.rd[37] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _25603_ (.A0(_01777_),
    .A1(_01773_),
    .S(_01683_),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _25604_ (.A0(mem_rdata[5]),
    .A1(mem_rdata[21]),
    .S(pcpi_rs1[1]),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _25605_ (.A0(_01774_),
    .A1(_01773_),
    .S(_00304_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _25606_ (.A0(_01768_),
    .A1(_01767_),
    .S(_01714_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _25607_ (.A0(_01770_),
    .A1(_01769_),
    .S(_01717_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _25608_ (.A0(\pcpi_mul.rd[4] ),
    .A1(\pcpi_mul.rd[36] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _25609_ (.A0(_01764_),
    .A1(_01760_),
    .S(_01683_),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _25610_ (.A0(mem_rdata[4]),
    .A1(mem_rdata[20]),
    .S(pcpi_rs1[1]),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _25611_ (.A0(_01761_),
    .A1(_01760_),
    .S(_00304_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _25612_ (.A0(_01755_),
    .A1(_01754_),
    .S(_01714_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _25613_ (.A0(_01757_),
    .A1(_01756_),
    .S(_01717_),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_1 _25614_ (.A0(\pcpi_mul.rd[3] ),
    .A1(\pcpi_mul.rd[35] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _25615_ (.A0(_01751_),
    .A1(_01747_),
    .S(_01683_),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _25616_ (.A0(mem_rdata[3]),
    .A1(mem_rdata[19]),
    .S(pcpi_rs1[1]),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _25617_ (.A0(_01748_),
    .A1(_01747_),
    .S(_00304_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _25618_ (.A0(_01742_),
    .A1(_01741_),
    .S(_01714_),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _25619_ (.A0(_01744_),
    .A1(_01743_),
    .S(_01717_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_1 _25620_ (.A0(\pcpi_mul.rd[2] ),
    .A1(\pcpi_mul.rd[34] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _25621_ (.A0(_01738_),
    .A1(_01734_),
    .S(_01683_),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _25622_ (.A0(mem_rdata[2]),
    .A1(mem_rdata[18]),
    .S(pcpi_rs1[1]),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _25623_ (.A0(_01735_),
    .A1(_01734_),
    .S(_00304_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_1 _25624_ (.A0(_01729_),
    .A1(_01728_),
    .S(_01714_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _25625_ (.A0(_01731_),
    .A1(_01730_),
    .S(_01717_),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_1 _25626_ (.A0(\pcpi_mul.rd[1] ),
    .A1(\pcpi_mul.rd[33] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _25627_ (.A0(_01725_),
    .A1(_01721_),
    .S(_01683_),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _25628_ (.A0(mem_rdata[1]),
    .A1(mem_rdata[17]),
    .S(pcpi_rs1[1]),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _25629_ (.A0(_01722_),
    .A1(_01721_),
    .S(_00304_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _25630_ (.A0(_01715_),
    .A1(_02559_),
    .S(_01714_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _25631_ (.A0(_01718_),
    .A1(_01716_),
    .S(_01717_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _25632_ (.A0(\pcpi_mul.rd[0] ),
    .A1(\pcpi_mul.rd[32] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _25633_ (.A0(_01711_),
    .A1(_01707_),
    .S(_01683_),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _25634_ (.A0(mem_rdata[0]),
    .A1(mem_rdata[16]),
    .S(pcpi_rs1[1]),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _25635_ (.A0(_01708_),
    .A1(_01707_),
    .S(_00304_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _25636_ (.A0(_01701_),
    .A1(_01696_),
    .S(_00311_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _25637_ (.A0(_01702_),
    .A1(_01696_),
    .S(\pcpi_mul.active[1] ),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _25638_ (.A0(_01696_),
    .A1(_01703_),
    .S(_00310_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _25639_ (.A0(_01693_),
    .A1(mem_wstrb[3]),
    .S(_00316_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _25640_ (.A0(_01690_),
    .A1(mem_wstrb[2]),
    .S(_00316_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _25641_ (.A0(_01687_),
    .A1(mem_wstrb[1]),
    .S(_00316_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _25642_ (.A0(_01684_),
    .A1(mem_wstrb[0]),
    .S(_00316_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _25643_ (.A0(\reg_next_pc[31] ),
    .A1(_01554_),
    .S(latched_store),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _25644_ (.A0(\reg_out[31] ),
    .A1(\alu_out_q[31] ),
    .S(latched_stalu),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _25645_ (.A0(\reg_next_pc[30] ),
    .A1(_01551_),
    .S(latched_store),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _25646_ (.A0(\reg_out[30] ),
    .A1(\alu_out_q[30] ),
    .S(latched_stalu),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _25647_ (.A0(\reg_next_pc[29] ),
    .A1(_01548_),
    .S(latched_store),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _25648_ (.A0(\reg_out[29] ),
    .A1(\alu_out_q[29] ),
    .S(latched_stalu),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _25649_ (.A0(\reg_next_pc[28] ),
    .A1(_01545_),
    .S(latched_store),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _25650_ (.A0(\reg_out[28] ),
    .A1(\alu_out_q[28] ),
    .S(latched_stalu),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _25651_ (.A0(\reg_next_pc[27] ),
    .A1(_01542_),
    .S(latched_store),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _25652_ (.A0(\reg_out[27] ),
    .A1(\alu_out_q[27] ),
    .S(latched_stalu),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _25653_ (.A0(\reg_next_pc[26] ),
    .A1(_01539_),
    .S(latched_store),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _25654_ (.A0(\reg_out[26] ),
    .A1(\alu_out_q[26] ),
    .S(latched_stalu),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _25655_ (.A0(\reg_next_pc[25] ),
    .A1(_01536_),
    .S(latched_store),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _25656_ (.A0(\reg_out[25] ),
    .A1(\alu_out_q[25] ),
    .S(latched_stalu),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _25657_ (.A0(\reg_next_pc[24] ),
    .A1(_01533_),
    .S(latched_store),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _25658_ (.A0(\reg_out[24] ),
    .A1(\alu_out_q[24] ),
    .S(latched_stalu),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _25659_ (.A0(\reg_next_pc[23] ),
    .A1(_01530_),
    .S(latched_store),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _25660_ (.A0(\reg_out[23] ),
    .A1(\alu_out_q[23] ),
    .S(latched_stalu),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _25661_ (.A0(\reg_next_pc[22] ),
    .A1(_01527_),
    .S(latched_store),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _25662_ (.A0(\reg_out[22] ),
    .A1(\alu_out_q[22] ),
    .S(latched_stalu),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _25663_ (.A0(\reg_next_pc[21] ),
    .A1(_01524_),
    .S(latched_store),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _25664_ (.A0(\reg_out[21] ),
    .A1(\alu_out_q[21] ),
    .S(latched_stalu),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _25665_ (.A0(\reg_next_pc[20] ),
    .A1(_01521_),
    .S(latched_store),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _25666_ (.A0(\reg_out[20] ),
    .A1(\alu_out_q[20] ),
    .S(latched_stalu),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _25667_ (.A0(\reg_next_pc[19] ),
    .A1(_01518_),
    .S(latched_store),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _25668_ (.A0(\reg_out[19] ),
    .A1(\alu_out_q[19] ),
    .S(latched_stalu),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _25669_ (.A0(\reg_next_pc[18] ),
    .A1(_01515_),
    .S(latched_store),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _25670_ (.A0(\reg_out[18] ),
    .A1(\alu_out_q[18] ),
    .S(latched_stalu),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _25671_ (.A0(\reg_next_pc[17] ),
    .A1(_01512_),
    .S(latched_store),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _25672_ (.A0(\reg_out[17] ),
    .A1(\alu_out_q[17] ),
    .S(latched_stalu),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _25673_ (.A0(\reg_next_pc[16] ),
    .A1(_01509_),
    .S(latched_store),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _25674_ (.A0(\reg_out[16] ),
    .A1(\alu_out_q[16] ),
    .S(latched_stalu),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _25675_ (.A0(\reg_next_pc[15] ),
    .A1(_01506_),
    .S(latched_store),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _25676_ (.A0(\reg_out[15] ),
    .A1(\alu_out_q[15] ),
    .S(latched_stalu),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _25677_ (.A0(\reg_next_pc[14] ),
    .A1(_01503_),
    .S(latched_store),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _25678_ (.A0(\reg_out[14] ),
    .A1(\alu_out_q[14] ),
    .S(latched_stalu),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _25679_ (.A0(\reg_next_pc[13] ),
    .A1(_01500_),
    .S(latched_store),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _25680_ (.A0(\reg_out[13] ),
    .A1(\alu_out_q[13] ),
    .S(latched_stalu),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _25681_ (.A0(\reg_next_pc[12] ),
    .A1(_01497_),
    .S(latched_store),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _25682_ (.A0(\reg_out[12] ),
    .A1(\alu_out_q[12] ),
    .S(latched_stalu),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _25683_ (.A0(\reg_next_pc[11] ),
    .A1(_01494_),
    .S(latched_store),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _25684_ (.A0(\reg_out[11] ),
    .A1(\alu_out_q[11] ),
    .S(latched_stalu),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _25685_ (.A0(\reg_next_pc[10] ),
    .A1(_01491_),
    .S(latched_store),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _25686_ (.A0(\reg_out[10] ),
    .A1(\alu_out_q[10] ),
    .S(latched_stalu),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _25687_ (.A0(\reg_next_pc[9] ),
    .A1(_01488_),
    .S(latched_store),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _25688_ (.A0(\reg_out[9] ),
    .A1(\alu_out_q[9] ),
    .S(latched_stalu),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _25689_ (.A0(\reg_next_pc[8] ),
    .A1(_01485_),
    .S(latched_store),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _25690_ (.A0(\reg_out[8] ),
    .A1(\alu_out_q[8] ),
    .S(latched_stalu),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _25691_ (.A0(\reg_next_pc[7] ),
    .A1(_01482_),
    .S(latched_store),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _25692_ (.A0(\reg_out[7] ),
    .A1(\alu_out_q[7] ),
    .S(latched_stalu),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _25693_ (.A0(\reg_next_pc[6] ),
    .A1(_01479_),
    .S(latched_store),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _25694_ (.A0(\reg_out[6] ),
    .A1(\alu_out_q[6] ),
    .S(latched_stalu),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _25695_ (.A0(\reg_next_pc[5] ),
    .A1(_01476_),
    .S(latched_store),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _25696_ (.A0(\reg_out[5] ),
    .A1(\alu_out_q[5] ),
    .S(latched_stalu),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _25697_ (.A0(_01474_),
    .A1(_01471_),
    .S(_00292_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _25698_ (.A0(\reg_next_pc[4] ),
    .A1(_01472_),
    .S(latched_store),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _25699_ (.A0(\reg_out[4] ),
    .A1(\alu_out_q[4] ),
    .S(latched_stalu),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _25700_ (.A0(\reg_next_pc[3] ),
    .A1(_01468_),
    .S(latched_store),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _25701_ (.A0(\reg_out[3] ),
    .A1(\alu_out_q[3] ),
    .S(latched_stalu),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _25702_ (.A0(\reg_next_pc[1] ),
    .A1(_01465_),
    .S(latched_store),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _25703_ (.A0(\reg_out[1] ),
    .A1(\alu_out_q[1] ),
    .S(latched_stalu),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _25704_ (.A0(_01301_),
    .A1(\timer[31] ),
    .S(_01208_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _25705_ (.A0(_01298_),
    .A1(\timer[30] ),
    .S(_01208_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _25706_ (.A0(_01295_),
    .A1(\timer[29] ),
    .S(_01208_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _25707_ (.A0(_01292_),
    .A1(\timer[28] ),
    .S(_01208_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _25708_ (.A0(_01289_),
    .A1(\timer[27] ),
    .S(_01208_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _25709_ (.A0(_01286_),
    .A1(\timer[26] ),
    .S(_01208_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _25710_ (.A0(_01283_),
    .A1(\timer[25] ),
    .S(_01208_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _25711_ (.A0(_01280_),
    .A1(\timer[24] ),
    .S(_01208_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _25712_ (.A0(_01277_),
    .A1(\timer[23] ),
    .S(_01208_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _25713_ (.A0(_01274_),
    .A1(\timer[22] ),
    .S(_01208_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _25714_ (.A0(_01271_),
    .A1(\timer[21] ),
    .S(_01208_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _25715_ (.A0(_01268_),
    .A1(\timer[20] ),
    .S(_01208_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _25716_ (.A0(_01265_),
    .A1(\timer[19] ),
    .S(_01208_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _25717_ (.A0(_01262_),
    .A1(\timer[18] ),
    .S(_01208_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _25718_ (.A0(_01259_),
    .A1(\timer[17] ),
    .S(_01208_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _25719_ (.A0(_01256_),
    .A1(\timer[16] ),
    .S(_01208_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _25720_ (.A0(_01253_),
    .A1(\timer[15] ),
    .S(_01208_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _25721_ (.A0(_01250_),
    .A1(\timer[14] ),
    .S(_01208_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _25722_ (.A0(_01247_),
    .A1(\timer[13] ),
    .S(_01208_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _25723_ (.A0(_01244_),
    .A1(\timer[12] ),
    .S(_01208_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _25724_ (.A0(_01241_),
    .A1(\timer[11] ),
    .S(_01208_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _25725_ (.A0(_01238_),
    .A1(\timer[10] ),
    .S(_01208_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _25726_ (.A0(_01235_),
    .A1(\timer[9] ),
    .S(_01208_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _25727_ (.A0(_01232_),
    .A1(\timer[8] ),
    .S(_01208_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _25728_ (.A0(_01229_),
    .A1(\timer[7] ),
    .S(_01208_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _25729_ (.A0(_01226_),
    .A1(\timer[6] ),
    .S(_01208_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _25730_ (.A0(_01223_),
    .A1(\timer[5] ),
    .S(_01208_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _25731_ (.A0(_01220_),
    .A1(\timer[4] ),
    .S(_01208_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _25732_ (.A0(_01217_),
    .A1(\timer[3] ),
    .S(_01208_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _25733_ (.A0(_01214_),
    .A1(\timer[2] ),
    .S(_01208_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _25734_ (.A0(_01211_),
    .A1(\timer[1] ),
    .S(_01208_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _25735_ (.A0(_01206_),
    .A1(_01201_),
    .S(_00368_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _25736_ (.A0(_01179_),
    .A1(_01174_),
    .S(_00368_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _25737_ (.A0(_01152_),
    .A1(_01147_),
    .S(_00368_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _25738_ (.A0(_01125_),
    .A1(_01120_),
    .S(_00368_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _25739_ (.A0(_01098_),
    .A1(_01093_),
    .S(_00368_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _25740_ (.A0(_01071_),
    .A1(_01066_),
    .S(_00368_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _25741_ (.A0(_01044_),
    .A1(_01039_),
    .S(_00368_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _25742_ (.A0(_01017_),
    .A1(_01012_),
    .S(_00368_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _25743_ (.A0(_00990_),
    .A1(_00985_),
    .S(_00368_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _25744_ (.A0(_00963_),
    .A1(_00958_),
    .S(_00368_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _25745_ (.A0(_00936_),
    .A1(_00931_),
    .S(_00368_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _25746_ (.A0(_00909_),
    .A1(_00904_),
    .S(_00368_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _25747_ (.A0(_00882_),
    .A1(_00877_),
    .S(_00368_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _25748_ (.A0(_00855_),
    .A1(_00850_),
    .S(_00368_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _25749_ (.A0(_00828_),
    .A1(_00823_),
    .S(_00368_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _25750_ (.A0(_00801_),
    .A1(_00796_),
    .S(_00368_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _25751_ (.A0(_00774_),
    .A1(_00769_),
    .S(_00368_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _25752_ (.A0(_00747_),
    .A1(_00742_),
    .S(_00368_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _25753_ (.A0(_00720_),
    .A1(_00715_),
    .S(_00368_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _25754_ (.A0(_00693_),
    .A1(_00688_),
    .S(_00368_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _25755_ (.A0(_00666_),
    .A1(_00661_),
    .S(_00368_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _25756_ (.A0(_00639_),
    .A1(_00634_),
    .S(_00368_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _25757_ (.A0(_00612_),
    .A1(_00607_),
    .S(_00368_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _25758_ (.A0(_00585_),
    .A1(_00580_),
    .S(_00368_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _25759_ (.A0(_00558_),
    .A1(_00553_),
    .S(_00368_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _25760_ (.A0(_00531_),
    .A1(_00526_),
    .S(_00368_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _25761_ (.A0(_00504_),
    .A1(_00499_),
    .S(_00368_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _25762_ (.A0(_00477_),
    .A1(_00472_),
    .S(_00368_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _25763_ (.A0(_00450_),
    .A1(_00445_),
    .S(_00368_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _25764_ (.A0(_00423_),
    .A1(_00418_),
    .S(_00368_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _25765_ (.A0(_00396_),
    .A1(_00391_),
    .S(_00368_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _25766_ (.A0(_00369_),
    .A1(_00365_),
    .S(_00368_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _25767_ (.A0(_00366_),
    .A1(_00367_),
    .S(\cpu_state[3] ),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _25768_ (.A0(\decoded_rs1[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(\cpu_state[3] ),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _25769_ (.A0(\decoded_rs1[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(\cpu_state[3] ),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _25770_ (.A0(\decoded_rs1[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(\cpu_state[3] ),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _25771_ (.A0(\decoded_rs1[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(\cpu_state[3] ),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _25772_ (.A0(_00349_),
    .A1(_00323_),
    .S(decoder_trigger),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _25773_ (.A0(_00350_),
    .A1(_00351_),
    .S(_00309_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _25774_ (.A0(_00352_),
    .A1(_00349_),
    .S(_00308_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _25775_ (.A0(_00355_),
    .A1(_00353_),
    .S(_00354_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _25776_ (.A0(_00337_),
    .A1(_00344_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _25777_ (.A0(_00345_),
    .A1(_00337_),
    .S(alu_wait),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _25778_ (.A0(_00342_),
    .A1(_00340_),
    .S(_00341_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _25779_ (.A0(_00338_),
    .A1(_00337_),
    .S(_00296_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _25780_ (.A0(\mem_rdata_q[12] ),
    .A1(_00334_),
    .S(\mem_rdata_q[13] ),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _25781_ (.A0(\cpu_state[1] ),
    .A1(_00302_),
    .S(\cpu_state[4] ),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _25782_ (.A0(_00322_),
    .A1(_00296_),
    .S(\cpu_state[6] ),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _25783_ (.A0(_00315_),
    .A1(alu_wait),
    .S(\cpu_state[4] ),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _25784_ (.A0(\mem_rdata_q[6] ),
    .A1(mem_rdata[6]),
    .S(mem_xfer),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _25785_ (.A0(\mem_rdata_q[5] ),
    .A1(mem_rdata[5]),
    .S(mem_xfer),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _25786_ (.A0(\mem_rdata_q[4] ),
    .A1(mem_rdata[4]),
    .S(mem_xfer),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _25787_ (.A0(\mem_rdata_q[3] ),
    .A1(mem_rdata[3]),
    .S(mem_xfer),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _25788_ (.A0(\mem_rdata_q[2] ),
    .A1(mem_rdata[2]),
    .S(mem_xfer),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _25789_ (.A0(\mem_rdata_q[1] ),
    .A1(mem_rdata[1]),
    .S(mem_xfer),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _25790_ (.A0(\mem_rdata_q[0] ),
    .A1(mem_rdata[0]),
    .S(mem_xfer),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _25791_ (.A0(\cpu_state[1] ),
    .A1(instr_retirq),
    .S(\cpu_state[2] ),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _25792_ (.A0(_00319_),
    .A1(\cpu_state[5] ),
    .S(_00296_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _25793_ (.A0(_00317_),
    .A1(\cpu_state[6] ),
    .S(_00296_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _25794_ (.A0(_00313_),
    .A1(_00312_),
    .S(_00307_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _25795_ (.A0(_00298_),
    .A1(_00299_),
    .S(_00289_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _25796_ (.A0(\reg_next_pc[2] ),
    .A1(_00293_),
    .S(latched_store),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _25797_ (.A0(\reg_out[2] ),
    .A1(\alu_out_q[2] ),
    .S(latched_stalu),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _25798_ (.A0(_00126_),
    .A1(_00122_),
    .S(mem_la_wdata[3]),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _25799_ (.A0(_00120_),
    .A1(_00116_),
    .S(mem_la_wdata[3]),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _25800_ (.A0(_00114_),
    .A1(_00110_),
    .S(mem_la_wdata[3]),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _25801_ (.A0(_00108_),
    .A1(_00104_),
    .S(mem_la_wdata[3]),
    .X(_02555_));
 sky130_fd_sc_hd__mux2_1 _25802_ (.A0(_00102_),
    .A1(_00095_),
    .S(mem_la_wdata[3]),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_1 _25803_ (.A0(_00092_),
    .A1(_00085_),
    .S(mem_la_wdata[3]),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_1 _25804_ (.A0(_00082_),
    .A1(_00068_),
    .S(mem_la_wdata[3]),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _25805_ (.A0(_00064_),
    .A1(_00050_),
    .S(mem_la_wdata[3]),
    .X(_02551_));
 sky130_fd_sc_hd__mux2_1 _25806_ (.A0(_01694_),
    .A1(_01695_),
    .S(_00290_),
    .X(_02541_));
 sky130_fd_sc_hd__mux2_1 _25807_ (.A0(_01691_),
    .A1(_01692_),
    .S(_00290_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _25808_ (.A0(_01688_),
    .A1(_01689_),
    .S(_00290_),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _25809_ (.A0(_01685_),
    .A1(_01686_),
    .S(_00290_),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _25810_ (.A0(_01679_),
    .A1(_01680_),
    .S(instr_jal),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _25811_ (.A0(_01682_),
    .A1(_02581_),
    .S(_00308_),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _25812_ (.A0(_01675_),
    .A1(_01676_),
    .S(instr_jal),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _25813_ (.A0(_01678_),
    .A1(_02580_),
    .S(_00308_),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _25814_ (.A0(_01671_),
    .A1(_01672_),
    .S(instr_jal),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _25815_ (.A0(_01674_),
    .A1(_02579_),
    .S(_00308_),
    .X(_02527_));
 sky130_fd_sc_hd__mux2_1 _25816_ (.A0(_01667_),
    .A1(_01668_),
    .S(instr_jal),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _25817_ (.A0(_01670_),
    .A1(_02578_),
    .S(_00308_),
    .X(_02526_));
 sky130_fd_sc_hd__mux2_1 _25818_ (.A0(_01663_),
    .A1(_01664_),
    .S(instr_jal),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _25819_ (.A0(_01666_),
    .A1(_02577_),
    .S(_00308_),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _25820_ (.A0(_01659_),
    .A1(_01660_),
    .S(instr_jal),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _25821_ (.A0(_01662_),
    .A1(_02576_),
    .S(_00308_),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _25822_ (.A0(_01655_),
    .A1(_01656_),
    .S(instr_jal),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _25823_ (.A0(_01658_),
    .A1(_02575_),
    .S(_00308_),
    .X(_02523_));
 sky130_fd_sc_hd__mux2_1 _25824_ (.A0(_01651_),
    .A1(_01652_),
    .S(instr_jal),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _25825_ (.A0(_01654_),
    .A1(_02574_),
    .S(_00308_),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _25826_ (.A0(_01647_),
    .A1(_01648_),
    .S(instr_jal),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _25827_ (.A0(_01650_),
    .A1(_02573_),
    .S(_00308_),
    .X(_02521_));
 sky130_fd_sc_hd__mux2_1 _25828_ (.A0(_01643_),
    .A1(_01644_),
    .S(instr_jal),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _25829_ (.A0(_01646_),
    .A1(_02572_),
    .S(_00308_),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _25830_ (.A0(_01639_),
    .A1(_01640_),
    .S(instr_jal),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _25831_ (.A0(_01642_),
    .A1(_02570_),
    .S(_00308_),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _25832_ (.A0(_01635_),
    .A1(_01636_),
    .S(instr_jal),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _25833_ (.A0(_01638_),
    .A1(_02569_),
    .S(_00308_),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _25834_ (.A0(_01631_),
    .A1(_01632_),
    .S(instr_jal),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _25835_ (.A0(_01634_),
    .A1(_02568_),
    .S(_00308_),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _25836_ (.A0(_01627_),
    .A1(_01628_),
    .S(instr_jal),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _25837_ (.A0(_01630_),
    .A1(_02567_),
    .S(_00308_),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _25838_ (.A0(_01623_),
    .A1(_01624_),
    .S(instr_jal),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _25839_ (.A0(_01626_),
    .A1(_02566_),
    .S(_00308_),
    .X(_02514_));
 sky130_fd_sc_hd__mux2_1 _25840_ (.A0(_01619_),
    .A1(_01620_),
    .S(instr_jal),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _25841_ (.A0(_01622_),
    .A1(_02565_),
    .S(_00308_),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _25842_ (.A0(_01615_),
    .A1(_01616_),
    .S(instr_jal),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _25843_ (.A0(_01618_),
    .A1(_02564_),
    .S(_00308_),
    .X(_02512_));
 sky130_fd_sc_hd__mux2_1 _25844_ (.A0(_01611_),
    .A1(_01612_),
    .S(instr_jal),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _25845_ (.A0(_01614_),
    .A1(_02563_),
    .S(_00308_),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _25846_ (.A0(_01607_),
    .A1(_01608_),
    .S(instr_jal),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _25847_ (.A0(_01610_),
    .A1(_02562_),
    .S(_00308_),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _25848_ (.A0(_01603_),
    .A1(_01604_),
    .S(instr_jal),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _25849_ (.A0(_01606_),
    .A1(_02561_),
    .S(_00308_),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _25850_ (.A0(_01599_),
    .A1(_01600_),
    .S(instr_jal),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _25851_ (.A0(_01602_),
    .A1(_02589_),
    .S(_00308_),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _25852_ (.A0(_01595_),
    .A1(_01596_),
    .S(instr_jal),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _25853_ (.A0(_01598_),
    .A1(_02588_),
    .S(_00308_),
    .X(_02507_));
 sky130_fd_sc_hd__mux2_1 _25854_ (.A0(_01591_),
    .A1(_01592_),
    .S(instr_jal),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _25855_ (.A0(_01594_),
    .A1(_02587_),
    .S(_00308_),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _25856_ (.A0(_01587_),
    .A1(_01588_),
    .S(instr_jal),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _25857_ (.A0(_01590_),
    .A1(_02586_),
    .S(_00308_),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _25858_ (.A0(_01583_),
    .A1(_01584_),
    .S(instr_jal),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _25859_ (.A0(_01586_),
    .A1(_02585_),
    .S(_00308_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _25860_ (.A0(_01579_),
    .A1(_01580_),
    .S(instr_jal),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _25861_ (.A0(_01582_),
    .A1(_02584_),
    .S(_00308_),
    .X(_02534_));
 sky130_fd_sc_hd__mux2_1 _25862_ (.A0(_01575_),
    .A1(_01576_),
    .S(instr_jal),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _25863_ (.A0(_01578_),
    .A1(_02583_),
    .S(_00308_),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _25864_ (.A0(_01571_),
    .A1(_01572_),
    .S(instr_jal),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _25865_ (.A0(_01574_),
    .A1(_02582_),
    .S(_00308_),
    .X(_02532_));
 sky130_fd_sc_hd__mux2_1 _25866_ (.A0(_01567_),
    .A1(_01568_),
    .S(instr_jal),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _25867_ (.A0(_01570_),
    .A1(_02571_),
    .S(_00308_),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _25868_ (.A0(_01561_),
    .A1(_01562_),
    .S(instr_jal),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _25869_ (.A0(_02560_),
    .A1(_01563_),
    .S(decoder_trigger),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _25870_ (.A0(_01564_),
    .A1(_01565_),
    .S(_00309_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _25871_ (.A0(_01566_),
    .A1(_02560_),
    .S(_00308_),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _25872_ (.A0(_02590_),
    .A1(_01557_),
    .S(instr_jal),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _25873_ (.A0(_02590_),
    .A1(_01558_),
    .S(decoder_trigger),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _25874_ (.A0(_01559_),
    .A1(_02590_),
    .S(_00309_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _25875_ (.A0(_01560_),
    .A1(_02590_),
    .S(_00308_),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _25876_ (.A0(\cpuregs_rs1[31] ),
    .A1(_01462_),
    .S(is_lui_auipc_jal),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _25877_ (.A0(_01464_),
    .A1(_01463_),
    .S(_00297_),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _25878_ (.A0(\cpuregs_rs1[30] ),
    .A1(_01459_),
    .S(is_lui_auipc_jal),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _25879_ (.A0(_01461_),
    .A1(_01460_),
    .S(_00297_),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _25880_ (.A0(\cpuregs_rs1[29] ),
    .A1(_01456_),
    .S(is_lui_auipc_jal),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _25881_ (.A0(_01458_),
    .A1(_01457_),
    .S(_00297_),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _25882_ (.A0(\cpuregs_rs1[28] ),
    .A1(_01453_),
    .S(is_lui_auipc_jal),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _25883_ (.A0(_01455_),
    .A1(_01454_),
    .S(_00297_),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _25884_ (.A0(\cpuregs_rs1[27] ),
    .A1(_01450_),
    .S(is_lui_auipc_jal),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _25885_ (.A0(_01452_),
    .A1(_01451_),
    .S(_00297_),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _25886_ (.A0(\cpuregs_rs1[26] ),
    .A1(_01447_),
    .S(is_lui_auipc_jal),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _25887_ (.A0(_01449_),
    .A1(_01448_),
    .S(_00297_),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _25888_ (.A0(\cpuregs_rs1[25] ),
    .A1(_01444_),
    .S(is_lui_auipc_jal),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _25889_ (.A0(_01446_),
    .A1(_01445_),
    .S(_00297_),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _25890_ (.A0(\cpuregs_rs1[24] ),
    .A1(_01441_),
    .S(is_lui_auipc_jal),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _25891_ (.A0(_01443_),
    .A1(_01442_),
    .S(_00297_),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _25892_ (.A0(\cpuregs_rs1[23] ),
    .A1(_01438_),
    .S(is_lui_auipc_jal),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _25893_ (.A0(_01440_),
    .A1(_01439_),
    .S(_00297_),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _25894_ (.A0(\cpuregs_rs1[22] ),
    .A1(_01435_),
    .S(is_lui_auipc_jal),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _25895_ (.A0(_01437_),
    .A1(_01436_),
    .S(_00297_),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _25896_ (.A0(\cpuregs_rs1[21] ),
    .A1(_01432_),
    .S(is_lui_auipc_jal),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _25897_ (.A0(_01434_),
    .A1(_01433_),
    .S(_00297_),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _25898_ (.A0(\cpuregs_rs1[20] ),
    .A1(_01429_),
    .S(is_lui_auipc_jal),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _25899_ (.A0(_01431_),
    .A1(_01430_),
    .S(_00297_),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _25900_ (.A0(\cpuregs_rs1[19] ),
    .A1(_01426_),
    .S(is_lui_auipc_jal),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _25901_ (.A0(_01428_),
    .A1(_01427_),
    .S(_00297_),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _25902_ (.A0(\cpuregs_rs1[18] ),
    .A1(_01423_),
    .S(is_lui_auipc_jal),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _25903_ (.A0(_01425_),
    .A1(_01424_),
    .S(_00297_),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _25904_ (.A0(\cpuregs_rs1[17] ),
    .A1(_01420_),
    .S(is_lui_auipc_jal),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _25905_ (.A0(_01422_),
    .A1(_01421_),
    .S(_00297_),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _25906_ (.A0(\cpuregs_rs1[16] ),
    .A1(_01417_),
    .S(is_lui_auipc_jal),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _25907_ (.A0(_01419_),
    .A1(_01418_),
    .S(_00297_),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _25908_ (.A0(\cpuregs_rs1[15] ),
    .A1(_01414_),
    .S(is_lui_auipc_jal),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _25909_ (.A0(_01416_),
    .A1(_01415_),
    .S(_00297_),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _25910_ (.A0(\cpuregs_rs1[14] ),
    .A1(_01411_),
    .S(is_lui_auipc_jal),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _25911_ (.A0(_01413_),
    .A1(_01412_),
    .S(_00297_),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _25912_ (.A0(\cpuregs_rs1[13] ),
    .A1(_01408_),
    .S(is_lui_auipc_jal),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _25913_ (.A0(_01410_),
    .A1(_01409_),
    .S(_00297_),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _25914_ (.A0(\cpuregs_rs1[12] ),
    .A1(_01405_),
    .S(is_lui_auipc_jal),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _25915_ (.A0(_01407_),
    .A1(_01406_),
    .S(_00297_),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _25916_ (.A0(\cpuregs_rs1[11] ),
    .A1(_01402_),
    .S(is_lui_auipc_jal),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _25917_ (.A0(_01404_),
    .A1(_01403_),
    .S(_00297_),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _25918_ (.A0(\cpuregs_rs1[10] ),
    .A1(_01399_),
    .S(is_lui_auipc_jal),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _25919_ (.A0(_01401_),
    .A1(_01400_),
    .S(_00297_),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _25920_ (.A0(\cpuregs_rs1[9] ),
    .A1(_01396_),
    .S(is_lui_auipc_jal),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _25921_ (.A0(_01398_),
    .A1(_01397_),
    .S(_00297_),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _25922_ (.A0(\cpuregs_rs1[8] ),
    .A1(_01393_),
    .S(is_lui_auipc_jal),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _25923_ (.A0(_01395_),
    .A1(_01394_),
    .S(_00297_),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_1 _25924_ (.A0(\cpuregs_rs1[7] ),
    .A1(_01390_),
    .S(is_lui_auipc_jal),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _25925_ (.A0(_01392_),
    .A1(_01391_),
    .S(_00297_),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _25926_ (.A0(\cpuregs_rs1[6] ),
    .A1(_01387_),
    .S(is_lui_auipc_jal),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _25927_ (.A0(_01389_),
    .A1(_01388_),
    .S(_00297_),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_1 _25928_ (.A0(\cpuregs_rs1[5] ),
    .A1(_01384_),
    .S(is_lui_auipc_jal),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _25929_ (.A0(_01386_),
    .A1(_01385_),
    .S(_00297_),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _25930_ (.A0(\cpuregs_rs1[4] ),
    .A1(_01381_),
    .S(is_lui_auipc_jal),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _25931_ (.A0(_01383_),
    .A1(_01382_),
    .S(_00297_),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _25932_ (.A0(\cpuregs_rs1[3] ),
    .A1(_01378_),
    .S(is_lui_auipc_jal),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _25933_ (.A0(_01380_),
    .A1(_01379_),
    .S(_00297_),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _25934_ (.A0(\cpuregs_rs1[2] ),
    .A1(_01375_),
    .S(is_lui_auipc_jal),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _25935_ (.A0(_01377_),
    .A1(_01376_),
    .S(_00297_),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _25936_ (.A0(\cpuregs_rs1[1] ),
    .A1(_01372_),
    .S(is_lui_auipc_jal),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _25937_ (.A0(_01374_),
    .A1(_01373_),
    .S(_00297_),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _25938_ (.A0(\cpuregs_rs1[0] ),
    .A1(_01369_),
    .S(is_lui_auipc_jal),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _25939_ (.A0(_01371_),
    .A1(_01370_),
    .S(_00297_),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _25940_ (.A0(_01367_),
    .A1(\decoded_imm[31] ),
    .S(_01304_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _25941_ (.A0(_01368_),
    .A1(\cpuregs_rs1[31] ),
    .S(\cpu_state[3] ),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _25942_ (.A0(_01365_),
    .A1(\decoded_imm[30] ),
    .S(_01304_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _25943_ (.A0(_01366_),
    .A1(\cpuregs_rs1[30] ),
    .S(\cpu_state[3] ),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _25944_ (.A0(_01363_),
    .A1(\decoded_imm[29] ),
    .S(_01304_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _25945_ (.A0(_01364_),
    .A1(\cpuregs_rs1[29] ),
    .S(\cpu_state[3] ),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _25946_ (.A0(_01361_),
    .A1(\decoded_imm[28] ),
    .S(_01304_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _25947_ (.A0(_01362_),
    .A1(\cpuregs_rs1[28] ),
    .S(\cpu_state[3] ),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _25948_ (.A0(_01359_),
    .A1(\decoded_imm[27] ),
    .S(_01304_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _25949_ (.A0(_01360_),
    .A1(\cpuregs_rs1[27] ),
    .S(\cpu_state[3] ),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _25950_ (.A0(_01357_),
    .A1(\decoded_imm[26] ),
    .S(_01304_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _25951_ (.A0(_01358_),
    .A1(\cpuregs_rs1[26] ),
    .S(\cpu_state[3] ),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _25952_ (.A0(_01355_),
    .A1(\decoded_imm[25] ),
    .S(_01304_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _25953_ (.A0(_01356_),
    .A1(\cpuregs_rs1[25] ),
    .S(\cpu_state[3] ),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _25954_ (.A0(_01353_),
    .A1(\decoded_imm[24] ),
    .S(_01304_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _25955_ (.A0(_01354_),
    .A1(\cpuregs_rs1[24] ),
    .S(\cpu_state[3] ),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _25956_ (.A0(_01351_),
    .A1(\decoded_imm[23] ),
    .S(_01304_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _25957_ (.A0(_01352_),
    .A1(\cpuregs_rs1[23] ),
    .S(\cpu_state[3] ),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _25958_ (.A0(_01349_),
    .A1(\decoded_imm[22] ),
    .S(_01304_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _25959_ (.A0(_01350_),
    .A1(\cpuregs_rs1[22] ),
    .S(\cpu_state[3] ),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _25960_ (.A0(_01347_),
    .A1(\decoded_imm[21] ),
    .S(_01304_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _25961_ (.A0(_01348_),
    .A1(\cpuregs_rs1[21] ),
    .S(\cpu_state[3] ),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _25962_ (.A0(_01345_),
    .A1(\decoded_imm[20] ),
    .S(_01304_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _25963_ (.A0(_01346_),
    .A1(\cpuregs_rs1[20] ),
    .S(\cpu_state[3] ),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _25964_ (.A0(_01343_),
    .A1(\decoded_imm[19] ),
    .S(_01304_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _25965_ (.A0(_01344_),
    .A1(\cpuregs_rs1[19] ),
    .S(\cpu_state[3] ),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _25966_ (.A0(_01341_),
    .A1(\decoded_imm[18] ),
    .S(_01304_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _25967_ (.A0(_01342_),
    .A1(\cpuregs_rs1[18] ),
    .S(\cpu_state[3] ),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _25968_ (.A0(_01339_),
    .A1(\decoded_imm[17] ),
    .S(_01304_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _25969_ (.A0(_01340_),
    .A1(\cpuregs_rs1[17] ),
    .S(\cpu_state[3] ),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _25970_ (.A0(_01337_),
    .A1(\decoded_imm[16] ),
    .S(_01304_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _25971_ (.A0(_01338_),
    .A1(\cpuregs_rs1[16] ),
    .S(\cpu_state[3] ),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _25972_ (.A0(_01335_),
    .A1(\decoded_imm[15] ),
    .S(_01304_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _25973_ (.A0(_01336_),
    .A1(\cpuregs_rs1[15] ),
    .S(\cpu_state[3] ),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _25974_ (.A0(_01333_),
    .A1(\decoded_imm[14] ),
    .S(_01304_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _25975_ (.A0(_01334_),
    .A1(\cpuregs_rs1[14] ),
    .S(\cpu_state[3] ),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _25976_ (.A0(_01331_),
    .A1(\decoded_imm[13] ),
    .S(_01304_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _25977_ (.A0(_01332_),
    .A1(\cpuregs_rs1[13] ),
    .S(\cpu_state[3] ),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _25978_ (.A0(_01329_),
    .A1(\decoded_imm[12] ),
    .S(_01304_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _25979_ (.A0(_01330_),
    .A1(\cpuregs_rs1[12] ),
    .S(\cpu_state[3] ),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _25980_ (.A0(_01327_),
    .A1(\decoded_imm[11] ),
    .S(_01304_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _25981_ (.A0(_01328_),
    .A1(\cpuregs_rs1[11] ),
    .S(\cpu_state[3] ),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _25982_ (.A0(_01325_),
    .A1(\decoded_imm[10] ),
    .S(_01304_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _25983_ (.A0(_01326_),
    .A1(\cpuregs_rs1[10] ),
    .S(\cpu_state[3] ),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _25984_ (.A0(_01323_),
    .A1(\decoded_imm[9] ),
    .S(_01304_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _25985_ (.A0(_01324_),
    .A1(\cpuregs_rs1[9] ),
    .S(\cpu_state[3] ),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _25986_ (.A0(_01321_),
    .A1(\decoded_imm[8] ),
    .S(_01304_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _25987_ (.A0(_01322_),
    .A1(\cpuregs_rs1[8] ),
    .S(\cpu_state[3] ),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _25988_ (.A0(_01319_),
    .A1(\decoded_imm[7] ),
    .S(_01304_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _25989_ (.A0(_01320_),
    .A1(\cpuregs_rs1[7] ),
    .S(\cpu_state[3] ),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _25990_ (.A0(_01317_),
    .A1(\decoded_imm[6] ),
    .S(_01304_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _25991_ (.A0(_01318_),
    .A1(\cpuregs_rs1[6] ),
    .S(\cpu_state[3] ),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _25992_ (.A0(_01315_),
    .A1(\decoded_imm[5] ),
    .S(_01304_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _25993_ (.A0(_01316_),
    .A1(\cpuregs_rs1[5] ),
    .S(\cpu_state[3] ),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _25994_ (.A0(\decoded_imm[4] ),
    .A1(\decoded_imm_uj[4] ),
    .S(is_slli_srli_srai),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _25995_ (.A0(_01313_),
    .A1(\decoded_imm[4] ),
    .S(_01304_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _25996_ (.A0(_01314_),
    .A1(\cpuregs_rs1[4] ),
    .S(\cpu_state[3] ),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _25997_ (.A0(\decoded_imm[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(is_slli_srli_srai),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _25998_ (.A0(_01311_),
    .A1(\decoded_imm[3] ),
    .S(_01304_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _25999_ (.A0(_01312_),
    .A1(\cpuregs_rs1[3] ),
    .S(\cpu_state[3] ),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _26000_ (.A0(\decoded_imm[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(is_slli_srli_srai),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _26001_ (.A0(_01309_),
    .A1(\decoded_imm[2] ),
    .S(_01304_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _26002_ (.A0(_01310_),
    .A1(\cpuregs_rs1[2] ),
    .S(\cpu_state[3] ),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _26003_ (.A0(\decoded_imm[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(is_slli_srli_srai),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _26004_ (.A0(_01307_),
    .A1(\decoded_imm[1] ),
    .S(_01304_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _26005_ (.A0(_01308_),
    .A1(\cpuregs_rs1[1] ),
    .S(\cpu_state[3] ),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _26006_ (.A0(\decoded_imm[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(is_slli_srli_srai),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _26007_ (.A0(_01305_),
    .A1(\decoded_imm[0] ),
    .S(_01304_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _26008_ (.A0(_01306_),
    .A1(\cpuregs_rs1[0] ),
    .S(\cpu_state[3] ),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _26009_ (.A0(_01302_),
    .A1(\cpuregs_rs1[31] ),
    .S(instr_timer),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _26010_ (.A0(_01302_),
    .A1(_01303_),
    .S(\cpu_state[2] ),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _26011_ (.A0(_01299_),
    .A1(\cpuregs_rs1[30] ),
    .S(instr_timer),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _26012_ (.A0(_01299_),
    .A1(_01300_),
    .S(\cpu_state[2] ),
    .X(_02434_));
 sky130_fd_sc_hd__mux2_1 _26013_ (.A0(_01296_),
    .A1(\cpuregs_rs1[29] ),
    .S(instr_timer),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _26014_ (.A0(_01296_),
    .A1(_01297_),
    .S(\cpu_state[2] ),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _26015_ (.A0(_01293_),
    .A1(\cpuregs_rs1[28] ),
    .S(instr_timer),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _26016_ (.A0(_01293_),
    .A1(_01294_),
    .S(\cpu_state[2] ),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _26017_ (.A0(_01290_),
    .A1(\cpuregs_rs1[27] ),
    .S(instr_timer),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _26018_ (.A0(_01290_),
    .A1(_01291_),
    .S(\cpu_state[2] ),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _26019_ (.A0(_01287_),
    .A1(\cpuregs_rs1[26] ),
    .S(instr_timer),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _26020_ (.A0(_01287_),
    .A1(_01288_),
    .S(\cpu_state[2] ),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _26021_ (.A0(_01284_),
    .A1(\cpuregs_rs1[25] ),
    .S(instr_timer),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _26022_ (.A0(_01284_),
    .A1(_01285_),
    .S(\cpu_state[2] ),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _26023_ (.A0(_01281_),
    .A1(\cpuregs_rs1[24] ),
    .S(instr_timer),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _26024_ (.A0(_01281_),
    .A1(_01282_),
    .S(\cpu_state[2] ),
    .X(_02427_));
 sky130_fd_sc_hd__mux2_1 _26025_ (.A0(_01278_),
    .A1(\cpuregs_rs1[23] ),
    .S(instr_timer),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _26026_ (.A0(_01278_),
    .A1(_01279_),
    .S(\cpu_state[2] ),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _26027_ (.A0(_01275_),
    .A1(\cpuregs_rs1[22] ),
    .S(instr_timer),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _26028_ (.A0(_01275_),
    .A1(_01276_),
    .S(\cpu_state[2] ),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _26029_ (.A0(_01272_),
    .A1(\cpuregs_rs1[21] ),
    .S(instr_timer),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _26030_ (.A0(_01272_),
    .A1(_01273_),
    .S(\cpu_state[2] ),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _26031_ (.A0(_01269_),
    .A1(\cpuregs_rs1[20] ),
    .S(instr_timer),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _26032_ (.A0(_01269_),
    .A1(_01270_),
    .S(\cpu_state[2] ),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _26033_ (.A0(_01266_),
    .A1(\cpuregs_rs1[19] ),
    .S(instr_timer),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _26034_ (.A0(_01266_),
    .A1(_01267_),
    .S(\cpu_state[2] ),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _26035_ (.A0(_01263_),
    .A1(\cpuregs_rs1[18] ),
    .S(instr_timer),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _26036_ (.A0(_01263_),
    .A1(_01264_),
    .S(\cpu_state[2] ),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _26037_ (.A0(_01260_),
    .A1(\cpuregs_rs1[17] ),
    .S(instr_timer),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _26038_ (.A0(_01260_),
    .A1(_01261_),
    .S(\cpu_state[2] ),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _26039_ (.A0(_01257_),
    .A1(\cpuregs_rs1[16] ),
    .S(instr_timer),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _26040_ (.A0(_01257_),
    .A1(_01258_),
    .S(\cpu_state[2] ),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _26041_ (.A0(_01254_),
    .A1(\cpuregs_rs1[15] ),
    .S(instr_timer),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _26042_ (.A0(_01254_),
    .A1(_01255_),
    .S(\cpu_state[2] ),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _26043_ (.A0(_01251_),
    .A1(\cpuregs_rs1[14] ),
    .S(instr_timer),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _26044_ (.A0(_01251_),
    .A1(_01252_),
    .S(\cpu_state[2] ),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _26045_ (.A0(_01248_),
    .A1(\cpuregs_rs1[13] ),
    .S(instr_timer),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _26046_ (.A0(_01248_),
    .A1(_01249_),
    .S(\cpu_state[2] ),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _26047_ (.A0(_01245_),
    .A1(\cpuregs_rs1[12] ),
    .S(instr_timer),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _26048_ (.A0(_01245_),
    .A1(_01246_),
    .S(\cpu_state[2] ),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _26049_ (.A0(_01242_),
    .A1(\cpuregs_rs1[11] ),
    .S(instr_timer),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _26050_ (.A0(_01242_),
    .A1(_01243_),
    .S(\cpu_state[2] ),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _26051_ (.A0(_01239_),
    .A1(\cpuregs_rs1[10] ),
    .S(instr_timer),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _26052_ (.A0(_01239_),
    .A1(_01240_),
    .S(\cpu_state[2] ),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _26053_ (.A0(_01236_),
    .A1(\cpuregs_rs1[9] ),
    .S(instr_timer),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _26054_ (.A0(_01236_),
    .A1(_01237_),
    .S(\cpu_state[2] ),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _26055_ (.A0(_01233_),
    .A1(\cpuregs_rs1[8] ),
    .S(instr_timer),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _26056_ (.A0(_01233_),
    .A1(_01234_),
    .S(\cpu_state[2] ),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _26057_ (.A0(_01230_),
    .A1(\cpuregs_rs1[7] ),
    .S(instr_timer),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _26058_ (.A0(_01230_),
    .A1(_01231_),
    .S(\cpu_state[2] ),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _26059_ (.A0(_01227_),
    .A1(\cpuregs_rs1[6] ),
    .S(instr_timer),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _26060_ (.A0(_01227_),
    .A1(_01228_),
    .S(\cpu_state[2] ),
    .X(_02439_));
 sky130_fd_sc_hd__mux2_1 _26061_ (.A0(_01224_),
    .A1(\cpuregs_rs1[5] ),
    .S(instr_timer),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _26062_ (.A0(_01224_),
    .A1(_01225_),
    .S(\cpu_state[2] ),
    .X(_02438_));
 sky130_fd_sc_hd__mux2_1 _26063_ (.A0(_01221_),
    .A1(\cpuregs_rs1[4] ),
    .S(instr_timer),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _26064_ (.A0(_01221_),
    .A1(_01222_),
    .S(\cpu_state[2] ),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _26065_ (.A0(_01218_),
    .A1(\cpuregs_rs1[3] ),
    .S(instr_timer),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _26066_ (.A0(_01218_),
    .A1(_01219_),
    .S(\cpu_state[2] ),
    .X(_02436_));
 sky130_fd_sc_hd__mux2_1 _26067_ (.A0(_01215_),
    .A1(\cpuregs_rs1[2] ),
    .S(instr_timer),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _26068_ (.A0(_01215_),
    .A1(_01216_),
    .S(\cpu_state[2] ),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_1 _26069_ (.A0(_01212_),
    .A1(\cpuregs_rs1[1] ),
    .S(instr_timer),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _26070_ (.A0(_01212_),
    .A1(_01213_),
    .S(\cpu_state[2] ),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _26071_ (.A0(_01209_),
    .A1(\cpuregs_rs1[0] ),
    .S(instr_timer),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _26072_ (.A0(_01209_),
    .A1(_01210_),
    .S(\cpu_state[2] ),
    .X(_02411_));
 sky130_fd_sc_hd__mux4_1 _26073_ (.A0(_01202_),
    .A1(_01203_),
    .A2(_01204_),
    .A3(_01205_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01206_));
 sky130_fd_sc_hd__mux4_1 _26074_ (.A0(_01181_),
    .A1(_01182_),
    .A2(_01183_),
    .A3(_01184_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01185_));
 sky130_fd_sc_hd__mux4_1 _26075_ (.A0(_01186_),
    .A1(_01187_),
    .A2(_01188_),
    .A3(_01189_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01190_));
 sky130_fd_sc_hd__mux4_1 _26076_ (.A0(_01191_),
    .A1(_01192_),
    .A2(_01193_),
    .A3(_01194_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01195_));
 sky130_fd_sc_hd__mux4_1 _26077_ (.A0(_01196_),
    .A1(_01197_),
    .A2(_01198_),
    .A3(_01199_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01200_));
 sky130_fd_sc_hd__mux4_1 _26078_ (.A0(_01185_),
    .A1(_01190_),
    .A2(_01195_),
    .A3(_01200_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01201_));
 sky130_fd_sc_hd__mux4_1 _26079_ (.A0(_01175_),
    .A1(_01176_),
    .A2(_01177_),
    .A3(_01178_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01179_));
 sky130_fd_sc_hd__mux4_1 _26080_ (.A0(_01154_),
    .A1(_01155_),
    .A2(_01156_),
    .A3(_01157_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01158_));
 sky130_fd_sc_hd__mux4_1 _26081_ (.A0(_01159_),
    .A1(_01160_),
    .A2(_01161_),
    .A3(_01162_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01163_));
 sky130_fd_sc_hd__mux4_1 _26082_ (.A0(_01164_),
    .A1(_01165_),
    .A2(_01166_),
    .A3(_01167_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01168_));
 sky130_fd_sc_hd__mux4_1 _26083_ (.A0(_01169_),
    .A1(_01170_),
    .A2(_01171_),
    .A3(_01172_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01173_));
 sky130_fd_sc_hd__mux4_1 _26084_ (.A0(_01158_),
    .A1(_01163_),
    .A2(_01168_),
    .A3(_01173_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01174_));
 sky130_fd_sc_hd__mux4_1 _26085_ (.A0(_01148_),
    .A1(_01149_),
    .A2(_01150_),
    .A3(_01151_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01152_));
 sky130_fd_sc_hd__mux4_1 _26086_ (.A0(_01127_),
    .A1(_01128_),
    .A2(_01129_),
    .A3(_01130_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01131_));
 sky130_fd_sc_hd__mux4_1 _26087_ (.A0(_01132_),
    .A1(_01133_),
    .A2(_01134_),
    .A3(_01135_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01136_));
 sky130_fd_sc_hd__mux4_1 _26088_ (.A0(_01137_),
    .A1(_01138_),
    .A2(_01139_),
    .A3(_01140_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01141_));
 sky130_fd_sc_hd__mux4_1 _26089_ (.A0(_01142_),
    .A1(_01143_),
    .A2(_01144_),
    .A3(_01145_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01146_));
 sky130_fd_sc_hd__mux4_1 _26090_ (.A0(_01131_),
    .A1(_01136_),
    .A2(_01141_),
    .A3(_01146_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01147_));
 sky130_fd_sc_hd__mux4_1 _26091_ (.A0(_01121_),
    .A1(_01122_),
    .A2(_01123_),
    .A3(_01124_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01125_));
 sky130_fd_sc_hd__mux4_1 _26092_ (.A0(_01100_),
    .A1(_01101_),
    .A2(_01102_),
    .A3(_01103_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01104_));
 sky130_fd_sc_hd__mux4_1 _26093_ (.A0(_01105_),
    .A1(_01106_),
    .A2(_01107_),
    .A3(_01108_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01109_));
 sky130_fd_sc_hd__mux4_1 _26094_ (.A0(_01110_),
    .A1(_01111_),
    .A2(_01112_),
    .A3(_01113_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01114_));
 sky130_fd_sc_hd__mux4_1 _26095_ (.A0(_01115_),
    .A1(_01116_),
    .A2(_01117_),
    .A3(_01118_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01119_));
 sky130_fd_sc_hd__mux4_1 _26096_ (.A0(_01104_),
    .A1(_01109_),
    .A2(_01114_),
    .A3(_01119_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01120_));
 sky130_fd_sc_hd__mux4_1 _26097_ (.A0(_01094_),
    .A1(_01095_),
    .A2(_01096_),
    .A3(_01097_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01098_));
 sky130_fd_sc_hd__mux4_1 _26098_ (.A0(_01073_),
    .A1(_01074_),
    .A2(_01075_),
    .A3(_01076_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01077_));
 sky130_fd_sc_hd__mux4_1 _26099_ (.A0(_01078_),
    .A1(_01079_),
    .A2(_01080_),
    .A3(_01081_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01082_));
 sky130_fd_sc_hd__mux4_1 _26100_ (.A0(_01083_),
    .A1(_01084_),
    .A2(_01085_),
    .A3(_01086_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01087_));
 sky130_fd_sc_hd__mux4_1 _26101_ (.A0(_01088_),
    .A1(_01089_),
    .A2(_01090_),
    .A3(_01091_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01092_));
 sky130_fd_sc_hd__mux4_1 _26102_ (.A0(_01077_),
    .A1(_01082_),
    .A2(_01087_),
    .A3(_01092_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01093_));
 sky130_fd_sc_hd__mux4_1 _26103_ (.A0(_01067_),
    .A1(_01068_),
    .A2(_01069_),
    .A3(_01070_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01071_));
 sky130_fd_sc_hd__mux4_1 _26104_ (.A0(_01046_),
    .A1(_01047_),
    .A2(_01048_),
    .A3(_01049_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01050_));
 sky130_fd_sc_hd__mux4_1 _26105_ (.A0(_01051_),
    .A1(_01052_),
    .A2(_01053_),
    .A3(_01054_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01055_));
 sky130_fd_sc_hd__mux4_1 _26106_ (.A0(_01056_),
    .A1(_01057_),
    .A2(_01058_),
    .A3(_01059_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01060_));
 sky130_fd_sc_hd__mux4_1 _26107_ (.A0(_01061_),
    .A1(_01062_),
    .A2(_01063_),
    .A3(_01064_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01065_));
 sky130_fd_sc_hd__mux4_1 _26108_ (.A0(_01050_),
    .A1(_01055_),
    .A2(_01060_),
    .A3(_01065_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01066_));
 sky130_fd_sc_hd__mux4_1 _26109_ (.A0(_01040_),
    .A1(_01041_),
    .A2(_01042_),
    .A3(_01043_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01044_));
 sky130_fd_sc_hd__mux4_1 _26110_ (.A0(_01019_),
    .A1(_01020_),
    .A2(_01021_),
    .A3(_01022_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01023_));
 sky130_fd_sc_hd__mux4_1 _26111_ (.A0(_01024_),
    .A1(_01025_),
    .A2(_01026_),
    .A3(_01027_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01028_));
 sky130_fd_sc_hd__mux4_1 _26112_ (.A0(_01029_),
    .A1(_01030_),
    .A2(_01031_),
    .A3(_01032_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01033_));
 sky130_fd_sc_hd__mux4_1 _26113_ (.A0(_01034_),
    .A1(_01035_),
    .A2(_01036_),
    .A3(_01037_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01038_));
 sky130_fd_sc_hd__mux4_1 _26114_ (.A0(_01023_),
    .A1(_01028_),
    .A2(_01033_),
    .A3(_01038_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01039_));
 sky130_fd_sc_hd__mux4_1 _26115_ (.A0(_01013_),
    .A1(_01014_),
    .A2(_01015_),
    .A3(_01016_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01017_));
 sky130_fd_sc_hd__mux4_1 _26116_ (.A0(_00992_),
    .A1(_00993_),
    .A2(_00994_),
    .A3(_00995_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00996_));
 sky130_fd_sc_hd__mux4_1 _26117_ (.A0(_00997_),
    .A1(_00998_),
    .A2(_00999_),
    .A3(_01000_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01001_));
 sky130_fd_sc_hd__mux4_1 _26118_ (.A0(_01002_),
    .A1(_01003_),
    .A2(_01004_),
    .A3(_01005_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01006_));
 sky130_fd_sc_hd__mux4_1 _26119_ (.A0(_01007_),
    .A1(_01008_),
    .A2(_01009_),
    .A3(_01010_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_01011_));
 sky130_fd_sc_hd__mux4_1 _26120_ (.A0(_00996_),
    .A1(_01001_),
    .A2(_01006_),
    .A3(_01011_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_01012_));
 sky130_fd_sc_hd__mux4_1 _26121_ (.A0(_00986_),
    .A1(_00987_),
    .A2(_00988_),
    .A3(_00989_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00990_));
 sky130_fd_sc_hd__mux4_1 _26122_ (.A0(_00965_),
    .A1(_00966_),
    .A2(_00967_),
    .A3(_00968_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00969_));
 sky130_fd_sc_hd__mux4_1 _26123_ (.A0(_00970_),
    .A1(_00971_),
    .A2(_00972_),
    .A3(_00973_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00974_));
 sky130_fd_sc_hd__mux4_1 _26124_ (.A0(_00975_),
    .A1(_00976_),
    .A2(_00977_),
    .A3(_00978_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00979_));
 sky130_fd_sc_hd__mux4_1 _26125_ (.A0(_00980_),
    .A1(_00981_),
    .A2(_00982_),
    .A3(_00983_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00984_));
 sky130_fd_sc_hd__mux4_1 _26126_ (.A0(_00969_),
    .A1(_00974_),
    .A2(_00979_),
    .A3(_00984_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00985_));
 sky130_fd_sc_hd__mux4_1 _26127_ (.A0(_00959_),
    .A1(_00960_),
    .A2(_00961_),
    .A3(_00962_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00963_));
 sky130_fd_sc_hd__mux4_1 _26128_ (.A0(_00938_),
    .A1(_00939_),
    .A2(_00940_),
    .A3(_00941_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00942_));
 sky130_fd_sc_hd__mux4_1 _26129_ (.A0(_00943_),
    .A1(_00944_),
    .A2(_00945_),
    .A3(_00946_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00947_));
 sky130_fd_sc_hd__mux4_1 _26130_ (.A0(_00948_),
    .A1(_00949_),
    .A2(_00950_),
    .A3(_00951_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00952_));
 sky130_fd_sc_hd__mux4_1 _26131_ (.A0(_00953_),
    .A1(_00954_),
    .A2(_00955_),
    .A3(_00956_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00957_));
 sky130_fd_sc_hd__mux4_1 _26132_ (.A0(_00942_),
    .A1(_00947_),
    .A2(_00952_),
    .A3(_00957_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00958_));
 sky130_fd_sc_hd__mux4_1 _26133_ (.A0(_00932_),
    .A1(_00933_),
    .A2(_00934_),
    .A3(_00935_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00936_));
 sky130_fd_sc_hd__mux4_1 _26134_ (.A0(_00911_),
    .A1(_00912_),
    .A2(_00913_),
    .A3(_00914_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00915_));
 sky130_fd_sc_hd__mux4_1 _26135_ (.A0(_00916_),
    .A1(_00917_),
    .A2(_00918_),
    .A3(_00919_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00920_));
 sky130_fd_sc_hd__mux4_1 _26136_ (.A0(_00921_),
    .A1(_00922_),
    .A2(_00923_),
    .A3(_00924_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00925_));
 sky130_fd_sc_hd__mux4_1 _26137_ (.A0(_00926_),
    .A1(_00927_),
    .A2(_00928_),
    .A3(_00929_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00930_));
 sky130_fd_sc_hd__mux4_1 _26138_ (.A0(_00915_),
    .A1(_00920_),
    .A2(_00925_),
    .A3(_00930_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00931_));
 sky130_fd_sc_hd__mux4_1 _26139_ (.A0(_00905_),
    .A1(_00906_),
    .A2(_00907_),
    .A3(_00908_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00909_));
 sky130_fd_sc_hd__mux4_1 _26140_ (.A0(_00884_),
    .A1(_00885_),
    .A2(_00886_),
    .A3(_00887_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00888_));
 sky130_fd_sc_hd__mux4_1 _26141_ (.A0(_00889_),
    .A1(_00890_),
    .A2(_00891_),
    .A3(_00892_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00893_));
 sky130_fd_sc_hd__mux4_1 _26142_ (.A0(_00894_),
    .A1(_00895_),
    .A2(_00896_),
    .A3(_00897_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00898_));
 sky130_fd_sc_hd__mux4_1 _26143_ (.A0(_00899_),
    .A1(_00900_),
    .A2(_00901_),
    .A3(_00902_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00903_));
 sky130_fd_sc_hd__mux4_1 _26144_ (.A0(_00888_),
    .A1(_00893_),
    .A2(_00898_),
    .A3(_00903_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00904_));
 sky130_fd_sc_hd__mux4_1 _26145_ (.A0(_00878_),
    .A1(_00879_),
    .A2(_00880_),
    .A3(_00881_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00882_));
 sky130_fd_sc_hd__mux4_1 _26146_ (.A0(_00857_),
    .A1(_00858_),
    .A2(_00859_),
    .A3(_00860_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00861_));
 sky130_fd_sc_hd__mux4_1 _26147_ (.A0(_00862_),
    .A1(_00863_),
    .A2(_00864_),
    .A3(_00865_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00866_));
 sky130_fd_sc_hd__mux4_1 _26148_ (.A0(_00867_),
    .A1(_00868_),
    .A2(_00869_),
    .A3(_00870_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00871_));
 sky130_fd_sc_hd__mux4_1 _26149_ (.A0(_00872_),
    .A1(_00873_),
    .A2(_00874_),
    .A3(_00875_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00876_));
 sky130_fd_sc_hd__mux4_1 _26150_ (.A0(_00861_),
    .A1(_00866_),
    .A2(_00871_),
    .A3(_00876_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00877_));
 sky130_fd_sc_hd__mux4_1 _26151_ (.A0(_00851_),
    .A1(_00852_),
    .A2(_00853_),
    .A3(_00854_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00855_));
 sky130_fd_sc_hd__mux4_1 _26152_ (.A0(_00830_),
    .A1(_00831_),
    .A2(_00832_),
    .A3(_00833_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00834_));
 sky130_fd_sc_hd__mux4_1 _26153_ (.A0(_00835_),
    .A1(_00836_),
    .A2(_00837_),
    .A3(_00838_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00839_));
 sky130_fd_sc_hd__mux4_1 _26154_ (.A0(_00840_),
    .A1(_00841_),
    .A2(_00842_),
    .A3(_00843_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00844_));
 sky130_fd_sc_hd__mux4_1 _26155_ (.A0(_00845_),
    .A1(_00846_),
    .A2(_00847_),
    .A3(_00848_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00849_));
 sky130_fd_sc_hd__mux4_1 _26156_ (.A0(_00834_),
    .A1(_00839_),
    .A2(_00844_),
    .A3(_00849_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00850_));
 sky130_fd_sc_hd__mux4_1 _26157_ (.A0(_00824_),
    .A1(_00825_),
    .A2(_00826_),
    .A3(_00827_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00828_));
 sky130_fd_sc_hd__mux4_1 _26158_ (.A0(_00803_),
    .A1(_00804_),
    .A2(_00805_),
    .A3(_00806_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00807_));
 sky130_fd_sc_hd__mux4_1 _26159_ (.A0(_00808_),
    .A1(_00809_),
    .A2(_00810_),
    .A3(_00811_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00812_));
 sky130_fd_sc_hd__mux4_1 _26160_ (.A0(_00813_),
    .A1(_00814_),
    .A2(_00815_),
    .A3(_00816_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00817_));
 sky130_fd_sc_hd__mux4_1 _26161_ (.A0(_00818_),
    .A1(_00819_),
    .A2(_00820_),
    .A3(_00821_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00822_));
 sky130_fd_sc_hd__mux4_1 _26162_ (.A0(_00807_),
    .A1(_00812_),
    .A2(_00817_),
    .A3(_00822_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00823_));
 sky130_fd_sc_hd__mux4_1 _26163_ (.A0(_00797_),
    .A1(_00798_),
    .A2(_00799_),
    .A3(_00800_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00801_));
 sky130_fd_sc_hd__mux4_1 _26164_ (.A0(_00776_),
    .A1(_00777_),
    .A2(_00778_),
    .A3(_00779_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00780_));
 sky130_fd_sc_hd__mux4_1 _26165_ (.A0(_00781_),
    .A1(_00782_),
    .A2(_00783_),
    .A3(_00784_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00785_));
 sky130_fd_sc_hd__mux4_1 _26166_ (.A0(_00786_),
    .A1(_00787_),
    .A2(_00788_),
    .A3(_00789_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00790_));
 sky130_fd_sc_hd__mux4_1 _26167_ (.A0(_00791_),
    .A1(_00792_),
    .A2(_00793_),
    .A3(_00794_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00795_));
 sky130_fd_sc_hd__mux4_1 _26168_ (.A0(_00780_),
    .A1(_00785_),
    .A2(_00790_),
    .A3(_00795_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00796_));
 sky130_fd_sc_hd__mux4_1 _26169_ (.A0(_00770_),
    .A1(_00771_),
    .A2(_00772_),
    .A3(_00773_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00774_));
 sky130_fd_sc_hd__mux4_1 _26170_ (.A0(_00749_),
    .A1(_00750_),
    .A2(_00751_),
    .A3(_00752_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00753_));
 sky130_fd_sc_hd__mux4_1 _26171_ (.A0(_00754_),
    .A1(_00755_),
    .A2(_00756_),
    .A3(_00757_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00758_));
 sky130_fd_sc_hd__mux4_1 _26172_ (.A0(_00759_),
    .A1(_00760_),
    .A2(_00761_),
    .A3(_00762_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00763_));
 sky130_fd_sc_hd__mux4_1 _26173_ (.A0(_00764_),
    .A1(_00765_),
    .A2(_00766_),
    .A3(_00767_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00768_));
 sky130_fd_sc_hd__mux4_1 _26174_ (.A0(_00753_),
    .A1(_00758_),
    .A2(_00763_),
    .A3(_00768_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00769_));
 sky130_fd_sc_hd__mux4_1 _26175_ (.A0(_00743_),
    .A1(_00744_),
    .A2(_00745_),
    .A3(_00746_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00747_));
 sky130_fd_sc_hd__mux4_1 _26176_ (.A0(_00722_),
    .A1(_00723_),
    .A2(_00724_),
    .A3(_00725_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00726_));
 sky130_fd_sc_hd__mux4_1 _26177_ (.A0(_00727_),
    .A1(_00728_),
    .A2(_00729_),
    .A3(_00730_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00731_));
 sky130_fd_sc_hd__mux4_1 _26178_ (.A0(_00732_),
    .A1(_00733_),
    .A2(_00734_),
    .A3(_00735_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00736_));
 sky130_fd_sc_hd__mux4_1 _26179_ (.A0(_00737_),
    .A1(_00738_),
    .A2(_00739_),
    .A3(_00740_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00741_));
 sky130_fd_sc_hd__mux4_1 _26180_ (.A0(_00726_),
    .A1(_00731_),
    .A2(_00736_),
    .A3(_00741_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00742_));
 sky130_fd_sc_hd__mux4_1 _26181_ (.A0(_00716_),
    .A1(_00717_),
    .A2(_00718_),
    .A3(_00719_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00720_));
 sky130_fd_sc_hd__mux4_1 _26182_ (.A0(_00695_),
    .A1(_00696_),
    .A2(_00697_),
    .A3(_00698_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00699_));
 sky130_fd_sc_hd__mux4_1 _26183_ (.A0(_00700_),
    .A1(_00701_),
    .A2(_00702_),
    .A3(_00703_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00704_));
 sky130_fd_sc_hd__mux4_1 _26184_ (.A0(_00705_),
    .A1(_00706_),
    .A2(_00707_),
    .A3(_00708_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00709_));
 sky130_fd_sc_hd__mux4_1 _26185_ (.A0(_00710_),
    .A1(_00711_),
    .A2(_00712_),
    .A3(_00713_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00714_));
 sky130_fd_sc_hd__mux4_1 _26186_ (.A0(_00699_),
    .A1(_00704_),
    .A2(_00709_),
    .A3(_00714_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00715_));
 sky130_fd_sc_hd__mux4_1 _26187_ (.A0(_00689_),
    .A1(_00690_),
    .A2(_00691_),
    .A3(_00692_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00693_));
 sky130_fd_sc_hd__mux4_1 _26188_ (.A0(_00668_),
    .A1(_00669_),
    .A2(_00670_),
    .A3(_00671_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00672_));
 sky130_fd_sc_hd__mux4_1 _26189_ (.A0(_00673_),
    .A1(_00674_),
    .A2(_00675_),
    .A3(_00676_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00677_));
 sky130_fd_sc_hd__mux4_1 _26190_ (.A0(_00678_),
    .A1(_00679_),
    .A2(_00680_),
    .A3(_00681_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00682_));
 sky130_fd_sc_hd__mux4_1 _26191_ (.A0(_00683_),
    .A1(_00684_),
    .A2(_00685_),
    .A3(_00686_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00687_));
 sky130_fd_sc_hd__mux4_1 _26192_ (.A0(_00672_),
    .A1(_00677_),
    .A2(_00682_),
    .A3(_00687_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00688_));
 sky130_fd_sc_hd__mux4_1 _26193_ (.A0(_00662_),
    .A1(_00663_),
    .A2(_00664_),
    .A3(_00665_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00666_));
 sky130_fd_sc_hd__mux4_1 _26194_ (.A0(_00641_),
    .A1(_00642_),
    .A2(_00643_),
    .A3(_00644_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00645_));
 sky130_fd_sc_hd__mux4_1 _26195_ (.A0(_00646_),
    .A1(_00647_),
    .A2(_00648_),
    .A3(_00649_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00650_));
 sky130_fd_sc_hd__mux4_1 _26196_ (.A0(_00651_),
    .A1(_00652_),
    .A2(_00653_),
    .A3(_00654_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00655_));
 sky130_fd_sc_hd__mux4_1 _26197_ (.A0(_00656_),
    .A1(_00657_),
    .A2(_00658_),
    .A3(_00659_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00660_));
 sky130_fd_sc_hd__mux4_1 _26198_ (.A0(_00645_),
    .A1(_00650_),
    .A2(_00655_),
    .A3(_00660_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00661_));
 sky130_fd_sc_hd__mux4_1 _26199_ (.A0(_00635_),
    .A1(_00636_),
    .A2(_00637_),
    .A3(_00638_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00639_));
 sky130_fd_sc_hd__mux4_1 _26200_ (.A0(_00614_),
    .A1(_00615_),
    .A2(_00616_),
    .A3(_00617_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00618_));
 sky130_fd_sc_hd__mux4_1 _26201_ (.A0(_00619_),
    .A1(_00620_),
    .A2(_00621_),
    .A3(_00622_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00623_));
 sky130_fd_sc_hd__mux4_1 _26202_ (.A0(_00624_),
    .A1(_00625_),
    .A2(_00626_),
    .A3(_00627_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00628_));
 sky130_fd_sc_hd__mux4_1 _26203_ (.A0(_00629_),
    .A1(_00630_),
    .A2(_00631_),
    .A3(_00632_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00633_));
 sky130_fd_sc_hd__mux4_1 _26204_ (.A0(_00618_),
    .A1(_00623_),
    .A2(_00628_),
    .A3(_00633_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00634_));
 sky130_fd_sc_hd__mux4_1 _26205_ (.A0(_00608_),
    .A1(_00609_),
    .A2(_00610_),
    .A3(_00611_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00612_));
 sky130_fd_sc_hd__mux4_1 _26206_ (.A0(_00587_),
    .A1(_00588_),
    .A2(_00589_),
    .A3(_00590_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00591_));
 sky130_fd_sc_hd__mux4_1 _26207_ (.A0(_00592_),
    .A1(_00593_),
    .A2(_00594_),
    .A3(_00595_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00596_));
 sky130_fd_sc_hd__mux4_1 _26208_ (.A0(_00597_),
    .A1(_00598_),
    .A2(_00599_),
    .A3(_00600_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00601_));
 sky130_fd_sc_hd__mux4_1 _26209_ (.A0(_00602_),
    .A1(_00603_),
    .A2(_00604_),
    .A3(_00605_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00606_));
 sky130_fd_sc_hd__mux4_1 _26210_ (.A0(_00591_),
    .A1(_00596_),
    .A2(_00601_),
    .A3(_00606_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00607_));
 sky130_fd_sc_hd__mux4_1 _26211_ (.A0(_00581_),
    .A1(_00582_),
    .A2(_00583_),
    .A3(_00584_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00585_));
 sky130_fd_sc_hd__mux4_1 _26212_ (.A0(_00560_),
    .A1(_00561_),
    .A2(_00562_),
    .A3(_00563_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00564_));
 sky130_fd_sc_hd__mux4_1 _26213_ (.A0(_00565_),
    .A1(_00566_),
    .A2(_00567_),
    .A3(_00568_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00569_));
 sky130_fd_sc_hd__mux4_1 _26214_ (.A0(_00570_),
    .A1(_00571_),
    .A2(_00572_),
    .A3(_00573_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00574_));
 sky130_fd_sc_hd__mux4_1 _26215_ (.A0(_00575_),
    .A1(_00576_),
    .A2(_00577_),
    .A3(_00578_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00579_));
 sky130_fd_sc_hd__mux4_1 _26216_ (.A0(_00564_),
    .A1(_00569_),
    .A2(_00574_),
    .A3(_00579_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00580_));
 sky130_fd_sc_hd__mux4_1 _26217_ (.A0(_00554_),
    .A1(_00555_),
    .A2(_00556_),
    .A3(_00557_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00558_));
 sky130_fd_sc_hd__mux4_1 _26218_ (.A0(_00533_),
    .A1(_00534_),
    .A2(_00535_),
    .A3(_00536_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00537_));
 sky130_fd_sc_hd__mux4_1 _26219_ (.A0(_00538_),
    .A1(_00539_),
    .A2(_00540_),
    .A3(_00541_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00542_));
 sky130_fd_sc_hd__mux4_1 _26220_ (.A0(_00543_),
    .A1(_00544_),
    .A2(_00545_),
    .A3(_00546_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00547_));
 sky130_fd_sc_hd__mux4_1 _26221_ (.A0(_00548_),
    .A1(_00549_),
    .A2(_00550_),
    .A3(_00551_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00552_));
 sky130_fd_sc_hd__mux4_1 _26222_ (.A0(_00537_),
    .A1(_00542_),
    .A2(_00547_),
    .A3(_00552_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00553_));
 sky130_fd_sc_hd__mux4_1 _26223_ (.A0(_00527_),
    .A1(_00528_),
    .A2(_00529_),
    .A3(_00530_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00531_));
 sky130_fd_sc_hd__mux4_1 _26224_ (.A0(_00506_),
    .A1(_00507_),
    .A2(_00508_),
    .A3(_00509_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00510_));
 sky130_fd_sc_hd__mux4_1 _26225_ (.A0(_00511_),
    .A1(_00512_),
    .A2(_00513_),
    .A3(_00514_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00515_));
 sky130_fd_sc_hd__mux4_1 _26226_ (.A0(_00516_),
    .A1(_00517_),
    .A2(_00518_),
    .A3(_00519_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00520_));
 sky130_fd_sc_hd__mux4_1 _26227_ (.A0(_00521_),
    .A1(_00522_),
    .A2(_00523_),
    .A3(_00524_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00525_));
 sky130_fd_sc_hd__mux4_1 _26228_ (.A0(_00510_),
    .A1(_00515_),
    .A2(_00520_),
    .A3(_00525_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00526_));
 sky130_fd_sc_hd__mux4_1 _26229_ (.A0(_00500_),
    .A1(_00501_),
    .A2(_00502_),
    .A3(_00503_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00504_));
 sky130_fd_sc_hd__mux4_1 _26230_ (.A0(_00479_),
    .A1(_00480_),
    .A2(_00481_),
    .A3(_00482_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00483_));
 sky130_fd_sc_hd__mux4_1 _26231_ (.A0(_00484_),
    .A1(_00485_),
    .A2(_00486_),
    .A3(_00487_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00488_));
 sky130_fd_sc_hd__mux4_1 _26232_ (.A0(_00489_),
    .A1(_00490_),
    .A2(_00491_),
    .A3(_00492_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00493_));
 sky130_fd_sc_hd__mux4_1 _26233_ (.A0(_00494_),
    .A1(_00495_),
    .A2(_00496_),
    .A3(_00497_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00498_));
 sky130_fd_sc_hd__mux4_1 _26234_ (.A0(_00483_),
    .A1(_00488_),
    .A2(_00493_),
    .A3(_00498_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00499_));
 sky130_fd_sc_hd__mux4_1 _26235_ (.A0(_00473_),
    .A1(_00474_),
    .A2(_00475_),
    .A3(_00476_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00477_));
 sky130_fd_sc_hd__mux4_1 _26236_ (.A0(_00452_),
    .A1(_00453_),
    .A2(_00454_),
    .A3(_00455_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00456_));
 sky130_fd_sc_hd__mux4_1 _26237_ (.A0(_00457_),
    .A1(_00458_),
    .A2(_00459_),
    .A3(_00460_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00461_));
 sky130_fd_sc_hd__mux4_1 _26238_ (.A0(_00462_),
    .A1(_00463_),
    .A2(_00464_),
    .A3(_00465_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00466_));
 sky130_fd_sc_hd__mux4_1 _26239_ (.A0(_00467_),
    .A1(_00468_),
    .A2(_00469_),
    .A3(_00470_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00471_));
 sky130_fd_sc_hd__mux4_1 _26240_ (.A0(_00456_),
    .A1(_00461_),
    .A2(_00466_),
    .A3(_00471_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00472_));
 sky130_fd_sc_hd__mux4_1 _26241_ (.A0(_00446_),
    .A1(_00447_),
    .A2(_00448_),
    .A3(_00449_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00450_));
 sky130_fd_sc_hd__mux4_1 _26242_ (.A0(_00425_),
    .A1(_00426_),
    .A2(_00427_),
    .A3(_00428_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00429_));
 sky130_fd_sc_hd__mux4_1 _26243_ (.A0(_00430_),
    .A1(_00431_),
    .A2(_00432_),
    .A3(_00433_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00434_));
 sky130_fd_sc_hd__mux4_1 _26244_ (.A0(_00435_),
    .A1(_00436_),
    .A2(_00437_),
    .A3(_00438_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00439_));
 sky130_fd_sc_hd__mux4_1 _26245_ (.A0(_00440_),
    .A1(_00441_),
    .A2(_00442_),
    .A3(_00443_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00444_));
 sky130_fd_sc_hd__mux4_1 _26246_ (.A0(_00429_),
    .A1(_00434_),
    .A2(_00439_),
    .A3(_00444_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00445_));
 sky130_fd_sc_hd__mux4_1 _26247_ (.A0(_00419_),
    .A1(_00420_),
    .A2(_00421_),
    .A3(_00422_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00423_));
 sky130_fd_sc_hd__mux4_1 _26248_ (.A0(_00398_),
    .A1(_00399_),
    .A2(_00400_),
    .A3(_00401_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00402_));
 sky130_fd_sc_hd__mux4_1 _26249_ (.A0(_00403_),
    .A1(_00404_),
    .A2(_00405_),
    .A3(_00406_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00407_));
 sky130_fd_sc_hd__mux4_1 _26250_ (.A0(_00408_),
    .A1(_00409_),
    .A2(_00410_),
    .A3(_00411_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00412_));
 sky130_fd_sc_hd__mux4_1 _26251_ (.A0(_00413_),
    .A1(_00414_),
    .A2(_00415_),
    .A3(_00416_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00417_));
 sky130_fd_sc_hd__mux4_1 _26252_ (.A0(_00402_),
    .A1(_00407_),
    .A2(_00412_),
    .A3(_00417_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00418_));
 sky130_fd_sc_hd__mux4_1 _26253_ (.A0(_00392_),
    .A1(_00393_),
    .A2(_00394_),
    .A3(_00395_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00396_));
 sky130_fd_sc_hd__mux4_1 _26254_ (.A0(_00371_),
    .A1(_00372_),
    .A2(_00373_),
    .A3(_00374_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00375_));
 sky130_fd_sc_hd__mux4_1 _26255_ (.A0(_00376_),
    .A1(_00377_),
    .A2(_00378_),
    .A3(_00379_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00380_));
 sky130_fd_sc_hd__mux4_1 _26256_ (.A0(_00381_),
    .A1(_00382_),
    .A2(_00383_),
    .A3(_00384_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00385_));
 sky130_fd_sc_hd__mux4_1 _26257_ (.A0(_00386_),
    .A1(_00387_),
    .A2(_00388_),
    .A3(_00389_),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00390_));
 sky130_fd_sc_hd__mux4_1 _26258_ (.A0(_00375_),
    .A1(_00380_),
    .A2(_00385_),
    .A3(_00390_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00391_));
 sky130_fd_sc_hd__mux4_1 _26259_ (.A0(\cpuregs[16][0] ),
    .A1(\cpuregs[17][0] ),
    .A2(\cpuregs[18][0] ),
    .A3(\cpuregs[19][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00369_));
 sky130_fd_sc_hd__mux4_1 _26260_ (.A0(\cpuregs[0][0] ),
    .A1(\cpuregs[1][0] ),
    .A2(\cpuregs[2][0] ),
    .A3(\cpuregs[3][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00359_));
 sky130_fd_sc_hd__mux4_1 _26261_ (.A0(\cpuregs[4][0] ),
    .A1(\cpuregs[5][0] ),
    .A2(\cpuregs[6][0] ),
    .A3(\cpuregs[7][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00361_));
 sky130_fd_sc_hd__mux4_1 _26262_ (.A0(\cpuregs[8][0] ),
    .A1(\cpuregs[9][0] ),
    .A2(\cpuregs[10][0] ),
    .A3(\cpuregs[11][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00363_));
 sky130_fd_sc_hd__mux4_1 _26263_ (.A0(\cpuregs[12][0] ),
    .A1(\cpuregs[13][0] ),
    .A2(\cpuregs[14][0] ),
    .A3(\cpuregs[15][0] ),
    .S0(_00357_),
    .S1(_00358_),
    .X(_00364_));
 sky130_fd_sc_hd__mux4_1 _26264_ (.A0(_00359_),
    .A1(_00361_),
    .A2(_00363_),
    .A3(_00364_),
    .S0(_00360_),
    .S1(_00362_),
    .X(_00365_));
 sky130_fd_sc_hd__mux4_1 _26265_ (.A0(_02581_),
    .A1(_01681_),
    .A2(_01679_),
    .A3(_02581_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01682_));
 sky130_fd_sc_hd__mux4_1 _26266_ (.A0(_02580_),
    .A1(_01677_),
    .A2(_01675_),
    .A3(_02580_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01678_));
 sky130_fd_sc_hd__mux4_1 _26267_ (.A0(_02579_),
    .A1(_01673_),
    .A2(_01671_),
    .A3(_02579_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01674_));
 sky130_fd_sc_hd__mux4_1 _26268_ (.A0(_02578_),
    .A1(_01669_),
    .A2(_01667_),
    .A3(_02578_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01670_));
 sky130_fd_sc_hd__mux4_1 _26269_ (.A0(_02577_),
    .A1(_01665_),
    .A2(_01663_),
    .A3(_02577_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01666_));
 sky130_fd_sc_hd__mux4_1 _26270_ (.A0(_02576_),
    .A1(_01661_),
    .A2(_01659_),
    .A3(_02576_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01662_));
 sky130_fd_sc_hd__mux4_1 _26271_ (.A0(_02575_),
    .A1(_01657_),
    .A2(_01655_),
    .A3(_02575_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01658_));
 sky130_fd_sc_hd__mux4_1 _26272_ (.A0(_02574_),
    .A1(_01653_),
    .A2(_01651_),
    .A3(_02574_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01654_));
 sky130_fd_sc_hd__mux4_1 _26273_ (.A0(_02573_),
    .A1(_01649_),
    .A2(_01647_),
    .A3(_02573_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01650_));
 sky130_fd_sc_hd__mux4_1 _26274_ (.A0(_02572_),
    .A1(_01645_),
    .A2(_01643_),
    .A3(_02572_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01646_));
 sky130_fd_sc_hd__mux4_1 _26275_ (.A0(_02570_),
    .A1(_01641_),
    .A2(_01639_),
    .A3(_02570_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01642_));
 sky130_fd_sc_hd__mux4_1 _26276_ (.A0(_02569_),
    .A1(_01637_),
    .A2(_01635_),
    .A3(_02569_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01638_));
 sky130_fd_sc_hd__mux4_1 _26277_ (.A0(_02568_),
    .A1(_01633_),
    .A2(_01631_),
    .A3(_02568_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01634_));
 sky130_fd_sc_hd__mux4_1 _26278_ (.A0(_02567_),
    .A1(_01629_),
    .A2(_01627_),
    .A3(_02567_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01630_));
 sky130_fd_sc_hd__mux4_1 _26279_ (.A0(_02566_),
    .A1(_01625_),
    .A2(_01623_),
    .A3(_02566_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01626_));
 sky130_fd_sc_hd__mux4_1 _26280_ (.A0(_02565_),
    .A1(_01621_),
    .A2(_01619_),
    .A3(_02565_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01622_));
 sky130_fd_sc_hd__mux4_1 _26281_ (.A0(_02564_),
    .A1(_01617_),
    .A2(_01615_),
    .A3(_02564_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01618_));
 sky130_fd_sc_hd__mux4_1 _26282_ (.A0(_02563_),
    .A1(_01613_),
    .A2(_01611_),
    .A3(_02563_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01614_));
 sky130_fd_sc_hd__mux4_1 _26283_ (.A0(_02562_),
    .A1(_01609_),
    .A2(_01607_),
    .A3(_02562_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01610_));
 sky130_fd_sc_hd__mux4_1 _26284_ (.A0(_02561_),
    .A1(_01605_),
    .A2(_01603_),
    .A3(_02561_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01606_));
 sky130_fd_sc_hd__mux4_1 _26285_ (.A0(_02589_),
    .A1(_01601_),
    .A2(_01599_),
    .A3(_02589_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01602_));
 sky130_fd_sc_hd__mux4_1 _26286_ (.A0(_02588_),
    .A1(_01597_),
    .A2(_01595_),
    .A3(_02588_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01598_));
 sky130_fd_sc_hd__mux4_1 _26287_ (.A0(_02587_),
    .A1(_01593_),
    .A2(_01591_),
    .A3(_02587_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01594_));
 sky130_fd_sc_hd__mux4_1 _26288_ (.A0(_02586_),
    .A1(_01589_),
    .A2(_01587_),
    .A3(_02586_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01590_));
 sky130_fd_sc_hd__mux4_1 _26289_ (.A0(_02585_),
    .A1(_01585_),
    .A2(_01583_),
    .A3(_02585_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01586_));
 sky130_fd_sc_hd__mux4_1 _26290_ (.A0(_02584_),
    .A1(_01581_),
    .A2(_01579_),
    .A3(_02584_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01582_));
 sky130_fd_sc_hd__mux4_1 _26291_ (.A0(_02583_),
    .A1(_01577_),
    .A2(_01575_),
    .A3(_02583_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01578_));
 sky130_fd_sc_hd__mux4_1 _26292_ (.A0(_02582_),
    .A1(_01573_),
    .A2(_01571_),
    .A3(_02582_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01574_));
 sky130_fd_sc_hd__mux4_1 _26293_ (.A0(_02571_),
    .A1(_01569_),
    .A2(_01567_),
    .A3(_02571_),
    .S0(_12946_),
    .S1(_00309_),
    .X(_01570_));
 sky130_fd_sc_hd__dfxtp_2 _26294_ (.CLK(clk),
    .D(_02687_),
    .Q(\alu_shl[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26295_ (.CLK(clk),
    .D(_02688_),
    .Q(\alu_shl[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26296_ (.CLK(clk),
    .D(_02689_),
    .Q(\alu_shl[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26297_ (.CLK(clk),
    .D(_02690_),
    .Q(\alu_shl[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26298_ (.CLK(clk),
    .D(_02691_),
    .Q(\alu_shl[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26299_ (.CLK(clk),
    .D(_02692_),
    .Q(\alu_shl[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26300_ (.CLK(clk),
    .D(_02693_),
    .Q(\alu_shl[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26301_ (.CLK(clk),
    .D(_02694_),
    .Q(\alu_shl[7] ));
 sky130_fd_sc_hd__dfxtp_2 _26302_ (.CLK(clk),
    .D(_02695_),
    .Q(\alu_shl[8] ));
 sky130_fd_sc_hd__dfxtp_2 _26303_ (.CLK(clk),
    .D(_02696_),
    .Q(\alu_shl[9] ));
 sky130_fd_sc_hd__dfxtp_2 _26304_ (.CLK(clk),
    .D(_02697_),
    .Q(\alu_shl[10] ));
 sky130_fd_sc_hd__dfxtp_2 _26305_ (.CLK(clk),
    .D(_02698_),
    .Q(\alu_shl[11] ));
 sky130_fd_sc_hd__dfxtp_2 _26306_ (.CLK(clk),
    .D(_02699_),
    .Q(\alu_shl[12] ));
 sky130_fd_sc_hd__dfxtp_2 _26307_ (.CLK(clk),
    .D(_02700_),
    .Q(\alu_shl[13] ));
 sky130_fd_sc_hd__dfxtp_2 _26308_ (.CLK(clk),
    .D(_02701_),
    .Q(\alu_shl[14] ));
 sky130_fd_sc_hd__dfxtp_2 _26309_ (.CLK(clk),
    .D(_02702_),
    .Q(\alu_shl[15] ));
 sky130_fd_sc_hd__dfxtp_2 _26310_ (.CLK(clk),
    .D(_02703_),
    .Q(alu_wait));
 sky130_fd_sc_hd__dfxtp_2 _26311_ (.CLK(clk),
    .D(_02704_),
    .Q(\latched_rd[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26312_ (.CLK(clk),
    .D(_02705_),
    .Q(\latched_rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26313_ (.CLK(clk),
    .D(_02706_),
    .Q(\latched_rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26314_ (.CLK(clk),
    .D(_02707_),
    .Q(\latched_rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26315_ (.CLK(clk),
    .D(_02708_),
    .Q(\decoded_imm[31] ));
 sky130_fd_sc_hd__dfxtp_2 _26316_ (.CLK(clk),
    .D(_02709_),
    .Q(\decoded_imm[30] ));
 sky130_fd_sc_hd__dfxtp_2 _26317_ (.CLK(clk),
    .D(_02710_),
    .Q(\decoded_imm[29] ));
 sky130_fd_sc_hd__dfxtp_2 _26318_ (.CLK(clk),
    .D(_02711_),
    .Q(\decoded_imm[28] ));
 sky130_fd_sc_hd__dfxtp_2 _26319_ (.CLK(clk),
    .D(_02712_),
    .Q(\decoded_imm[27] ));
 sky130_fd_sc_hd__dfxtp_2 _26320_ (.CLK(clk),
    .D(_02713_),
    .Q(\decoded_imm[26] ));
 sky130_fd_sc_hd__dfxtp_2 _26321_ (.CLK(clk),
    .D(_02714_),
    .Q(\decoded_imm[25] ));
 sky130_fd_sc_hd__dfxtp_2 _26322_ (.CLK(clk),
    .D(_02715_),
    .Q(\decoded_imm[24] ));
 sky130_fd_sc_hd__dfxtp_2 _26323_ (.CLK(clk),
    .D(_02716_),
    .Q(\decoded_imm[23] ));
 sky130_fd_sc_hd__dfxtp_2 _26324_ (.CLK(clk),
    .D(_02717_),
    .Q(\decoded_imm[22] ));
 sky130_fd_sc_hd__dfxtp_2 _26325_ (.CLK(clk),
    .D(_02718_),
    .Q(\decoded_imm[21] ));
 sky130_fd_sc_hd__dfxtp_2 _26326_ (.CLK(clk),
    .D(_02719_),
    .Q(\decoded_imm[20] ));
 sky130_fd_sc_hd__dfxtp_2 _26327_ (.CLK(clk),
    .D(_02720_),
    .Q(\decoded_imm[19] ));
 sky130_fd_sc_hd__dfxtp_2 _26328_ (.CLK(clk),
    .D(_02721_),
    .Q(\decoded_imm[18] ));
 sky130_fd_sc_hd__dfxtp_2 _26329_ (.CLK(clk),
    .D(_02722_),
    .Q(\decoded_imm[17] ));
 sky130_fd_sc_hd__dfxtp_2 _26330_ (.CLK(clk),
    .D(_02723_),
    .Q(\decoded_imm[16] ));
 sky130_fd_sc_hd__dfxtp_2 _26331_ (.CLK(clk),
    .D(_02724_),
    .Q(\decoded_imm[15] ));
 sky130_fd_sc_hd__dfxtp_2 _26332_ (.CLK(clk),
    .D(_02725_),
    .Q(\decoded_imm[14] ));
 sky130_fd_sc_hd__dfxtp_2 _26333_ (.CLK(clk),
    .D(_02726_),
    .Q(\decoded_imm[13] ));
 sky130_fd_sc_hd__dfxtp_2 _26334_ (.CLK(clk),
    .D(_02727_),
    .Q(\decoded_imm[12] ));
 sky130_fd_sc_hd__dfxtp_2 _26335_ (.CLK(clk),
    .D(_02728_),
    .Q(\decoded_imm[11] ));
 sky130_fd_sc_hd__dfxtp_2 _26336_ (.CLK(clk),
    .D(_02729_),
    .Q(\decoded_imm[10] ));
 sky130_fd_sc_hd__dfxtp_2 _26337_ (.CLK(clk),
    .D(_02730_),
    .Q(\decoded_imm[9] ));
 sky130_fd_sc_hd__dfxtp_2 _26338_ (.CLK(clk),
    .D(_02731_),
    .Q(\decoded_imm[8] ));
 sky130_fd_sc_hd__dfxtp_2 _26339_ (.CLK(clk),
    .D(_02732_),
    .Q(\decoded_imm[7] ));
 sky130_fd_sc_hd__dfxtp_2 _26340_ (.CLK(clk),
    .D(_02733_),
    .Q(\decoded_imm[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26341_ (.CLK(clk),
    .D(_02734_),
    .Q(\decoded_imm[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26342_ (.CLK(clk),
    .D(_02735_),
    .Q(\decoded_imm[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26343_ (.CLK(clk),
    .D(_02736_),
    .Q(\decoded_imm[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26344_ (.CLK(clk),
    .D(_02737_),
    .Q(\decoded_imm[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26345_ (.CLK(clk),
    .D(_02738_),
    .Q(\decoded_imm[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26346_ (.CLK(clk),
    .D(_02739_),
    .Q(\irq_pending[31] ));
 sky130_fd_sc_hd__dfxtp_2 _26347_ (.CLK(clk),
    .D(_02740_),
    .Q(\irq_pending[30] ));
 sky130_fd_sc_hd__dfxtp_2 _26348_ (.CLK(clk),
    .D(_02741_),
    .Q(\irq_pending[29] ));
 sky130_fd_sc_hd__dfxtp_2 _26349_ (.CLK(clk),
    .D(_02742_),
    .Q(\irq_pending[28] ));
 sky130_fd_sc_hd__dfxtp_2 _26350_ (.CLK(clk),
    .D(_02743_),
    .Q(\irq_pending[27] ));
 sky130_fd_sc_hd__dfxtp_2 _26351_ (.CLK(clk),
    .D(_02744_),
    .Q(\irq_pending[26] ));
 sky130_fd_sc_hd__dfxtp_2 _26352_ (.CLK(clk),
    .D(_02745_),
    .Q(\irq_pending[25] ));
 sky130_fd_sc_hd__dfxtp_2 _26353_ (.CLK(clk),
    .D(_02746_),
    .Q(\irq_pending[24] ));
 sky130_fd_sc_hd__dfxtp_2 _26354_ (.CLK(clk),
    .D(_02747_),
    .Q(\irq_pending[23] ));
 sky130_fd_sc_hd__dfxtp_2 _26355_ (.CLK(clk),
    .D(_02748_),
    .Q(\irq_pending[22] ));
 sky130_fd_sc_hd__dfxtp_2 _26356_ (.CLK(clk),
    .D(_02749_),
    .Q(\irq_pending[21] ));
 sky130_fd_sc_hd__dfxtp_2 _26357_ (.CLK(clk),
    .D(_02750_),
    .Q(\irq_pending[20] ));
 sky130_fd_sc_hd__dfxtp_2 _26358_ (.CLK(clk),
    .D(_02751_),
    .Q(\irq_pending[19] ));
 sky130_fd_sc_hd__dfxtp_2 _26359_ (.CLK(clk),
    .D(_02752_),
    .Q(\irq_pending[18] ));
 sky130_fd_sc_hd__dfxtp_2 _26360_ (.CLK(clk),
    .D(_02753_),
    .Q(\irq_pending[17] ));
 sky130_fd_sc_hd__dfxtp_2 _26361_ (.CLK(clk),
    .D(_02754_),
    .Q(\irq_pending[16] ));
 sky130_fd_sc_hd__dfxtp_2 _26362_ (.CLK(clk),
    .D(_02755_),
    .Q(\irq_pending[15] ));
 sky130_fd_sc_hd__dfxtp_2 _26363_ (.CLK(clk),
    .D(_02756_),
    .Q(\irq_pending[14] ));
 sky130_fd_sc_hd__dfxtp_2 _26364_ (.CLK(clk),
    .D(_02757_),
    .Q(\irq_pending[13] ));
 sky130_fd_sc_hd__dfxtp_2 _26365_ (.CLK(clk),
    .D(_02758_),
    .Q(\irq_pending[12] ));
 sky130_fd_sc_hd__dfxtp_2 _26366_ (.CLK(clk),
    .D(_02759_),
    .Q(\irq_pending[11] ));
 sky130_fd_sc_hd__dfxtp_2 _26367_ (.CLK(clk),
    .D(_02760_),
    .Q(\irq_pending[10] ));
 sky130_fd_sc_hd__dfxtp_2 _26368_ (.CLK(clk),
    .D(_02761_),
    .Q(\irq_pending[9] ));
 sky130_fd_sc_hd__dfxtp_2 _26369_ (.CLK(clk),
    .D(_02762_),
    .Q(\irq_pending[8] ));
 sky130_fd_sc_hd__dfxtp_2 _26370_ (.CLK(clk),
    .D(_02763_),
    .Q(\irq_pending[7] ));
 sky130_fd_sc_hd__dfxtp_2 _26371_ (.CLK(clk),
    .D(_02764_),
    .Q(\irq_pending[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26372_ (.CLK(clk),
    .D(_02765_),
    .Q(\irq_pending[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26373_ (.CLK(clk),
    .D(_02766_),
    .Q(\irq_pending[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26374_ (.CLK(clk),
    .D(_02767_),
    .Q(\irq_pending[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26375_ (.CLK(clk),
    .D(_02768_),
    .Q(\irq_pending[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26376_ (.CLK(clk),
    .D(_02769_),
    .Q(\irq_pending[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26377_ (.CLK(clk),
    .D(_02770_),
    .Q(\reg_next_pc[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26378_ (.CLK(clk),
    .D(_00045_),
    .Q(\mem_wordsize[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26379_ (.CLK(clk),
    .D(_00046_),
    .Q(\mem_wordsize[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26380_ (.CLK(clk),
    .D(_00047_),
    .Q(\mem_wordsize[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26381_ (.CLK(clk),
    .D(_12948_),
    .Q(\reg_out[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26382_ (.CLK(clk),
    .D(_12959_),
    .Q(\reg_out[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26383_ (.CLK(clk),
    .D(_12970_),
    .Q(\reg_out[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26384_ (.CLK(clk),
    .D(_12973_),
    .Q(\reg_out[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26385_ (.CLK(clk),
    .D(_12974_),
    .Q(\reg_out[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26386_ (.CLK(clk),
    .D(_12975_),
    .Q(\reg_out[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26387_ (.CLK(clk),
    .D(_12976_),
    .Q(\reg_out[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26388_ (.CLK(clk),
    .D(_12977_),
    .Q(\reg_out[7] ));
 sky130_fd_sc_hd__dfxtp_2 _26389_ (.CLK(clk),
    .D(_12978_),
    .Q(\reg_out[8] ));
 sky130_fd_sc_hd__dfxtp_2 _26390_ (.CLK(clk),
    .D(_12979_),
    .Q(\reg_out[9] ));
 sky130_fd_sc_hd__dfxtp_2 _26391_ (.CLK(clk),
    .D(_12949_),
    .Q(\reg_out[10] ));
 sky130_fd_sc_hd__dfxtp_2 _26392_ (.CLK(clk),
    .D(_12950_),
    .Q(\reg_out[11] ));
 sky130_fd_sc_hd__dfxtp_2 _26393_ (.CLK(clk),
    .D(_12951_),
    .Q(\reg_out[12] ));
 sky130_fd_sc_hd__dfxtp_2 _26394_ (.CLK(clk),
    .D(_12952_),
    .Q(\reg_out[13] ));
 sky130_fd_sc_hd__dfxtp_2 _26395_ (.CLK(clk),
    .D(_12953_),
    .Q(\reg_out[14] ));
 sky130_fd_sc_hd__dfxtp_2 _26396_ (.CLK(clk),
    .D(_12954_),
    .Q(\reg_out[15] ));
 sky130_fd_sc_hd__dfxtp_2 _26397_ (.CLK(clk),
    .D(_12955_),
    .Q(\reg_out[16] ));
 sky130_fd_sc_hd__dfxtp_2 _26398_ (.CLK(clk),
    .D(_12956_),
    .Q(\reg_out[17] ));
 sky130_fd_sc_hd__dfxtp_2 _26399_ (.CLK(clk),
    .D(_12957_),
    .Q(\reg_out[18] ));
 sky130_fd_sc_hd__dfxtp_2 _26400_ (.CLK(clk),
    .D(_12958_),
    .Q(\reg_out[19] ));
 sky130_fd_sc_hd__dfxtp_2 _26401_ (.CLK(clk),
    .D(_12960_),
    .Q(\reg_out[20] ));
 sky130_fd_sc_hd__dfxtp_2 _26402_ (.CLK(clk),
    .D(_12961_),
    .Q(\reg_out[21] ));
 sky130_fd_sc_hd__dfxtp_2 _26403_ (.CLK(clk),
    .D(_12962_),
    .Q(\reg_out[22] ));
 sky130_fd_sc_hd__dfxtp_2 _26404_ (.CLK(clk),
    .D(_12963_),
    .Q(\reg_out[23] ));
 sky130_fd_sc_hd__dfxtp_2 _26405_ (.CLK(clk),
    .D(_12964_),
    .Q(\reg_out[24] ));
 sky130_fd_sc_hd__dfxtp_2 _26406_ (.CLK(clk),
    .D(_12965_),
    .Q(\reg_out[25] ));
 sky130_fd_sc_hd__dfxtp_2 _26407_ (.CLK(clk),
    .D(_12966_),
    .Q(\reg_out[26] ));
 sky130_fd_sc_hd__dfxtp_2 _26408_ (.CLK(clk),
    .D(_12967_),
    .Q(\reg_out[27] ));
 sky130_fd_sc_hd__dfxtp_2 _26409_ (.CLK(clk),
    .D(_12968_),
    .Q(\reg_out[28] ));
 sky130_fd_sc_hd__dfxtp_2 _26410_ (.CLK(clk),
    .D(_12969_),
    .Q(\reg_out[29] ));
 sky130_fd_sc_hd__dfxtp_2 _26411_ (.CLK(clk),
    .D(_12971_),
    .Q(\reg_out[30] ));
 sky130_fd_sc_hd__dfxtp_2 _26412_ (.CLK(clk),
    .D(_12972_),
    .Q(\reg_out[31] ));
 sky130_fd_sc_hd__dfxtp_2 _26413_ (.CLK(clk),
    .D(_00004_),
    .Q(\irq_pending[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26414_ (.CLK(clk),
    .D(_00003_),
    .Q(decoder_trigger));
 sky130_fd_sc_hd__dfxtp_2 _26415_ (.CLK(clk),
    .D(\alu_out[0] ),
    .Q(\alu_out_q[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26416_ (.CLK(clk),
    .D(\alu_out[1] ),
    .Q(\alu_out_q[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26417_ (.CLK(clk),
    .D(\alu_out[2] ),
    .Q(\alu_out_q[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26418_ (.CLK(clk),
    .D(\alu_out[3] ),
    .Q(\alu_out_q[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26419_ (.CLK(clk),
    .D(\alu_out[4] ),
    .Q(\alu_out_q[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26420_ (.CLK(clk),
    .D(\alu_out[5] ),
    .Q(\alu_out_q[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26421_ (.CLK(clk),
    .D(\alu_out[6] ),
    .Q(\alu_out_q[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26422_ (.CLK(clk),
    .D(\alu_out[7] ),
    .Q(\alu_out_q[7] ));
 sky130_fd_sc_hd__dfxtp_2 _26423_ (.CLK(clk),
    .D(\alu_out[8] ),
    .Q(\alu_out_q[8] ));
 sky130_fd_sc_hd__dfxtp_2 _26424_ (.CLK(clk),
    .D(\alu_out[9] ),
    .Q(\alu_out_q[9] ));
 sky130_fd_sc_hd__dfxtp_2 _26425_ (.CLK(clk),
    .D(\alu_out[10] ),
    .Q(\alu_out_q[10] ));
 sky130_fd_sc_hd__dfxtp_2 _26426_ (.CLK(clk),
    .D(\alu_out[11] ),
    .Q(\alu_out_q[11] ));
 sky130_fd_sc_hd__dfxtp_2 _26427_ (.CLK(clk),
    .D(\alu_out[12] ),
    .Q(\alu_out_q[12] ));
 sky130_fd_sc_hd__dfxtp_2 _26428_ (.CLK(clk),
    .D(\alu_out[13] ),
    .Q(\alu_out_q[13] ));
 sky130_fd_sc_hd__dfxtp_2 _26429_ (.CLK(clk),
    .D(\alu_out[14] ),
    .Q(\alu_out_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _26430_ (.CLK(clk),
    .D(\alu_out[15] ),
    .Q(\alu_out_q[15] ));
 sky130_fd_sc_hd__dfxtp_2 _26431_ (.CLK(clk),
    .D(\alu_out[16] ),
    .Q(\alu_out_q[16] ));
 sky130_fd_sc_hd__dfxtp_2 _26432_ (.CLK(clk),
    .D(\alu_out[17] ),
    .Q(\alu_out_q[17] ));
 sky130_fd_sc_hd__dfxtp_2 _26433_ (.CLK(clk),
    .D(\alu_out[18] ),
    .Q(\alu_out_q[18] ));
 sky130_fd_sc_hd__dfxtp_2 _26434_ (.CLK(clk),
    .D(\alu_out[19] ),
    .Q(\alu_out_q[19] ));
 sky130_fd_sc_hd__dfxtp_2 _26435_ (.CLK(clk),
    .D(\alu_out[20] ),
    .Q(\alu_out_q[20] ));
 sky130_fd_sc_hd__dfxtp_2 _26436_ (.CLK(clk),
    .D(\alu_out[21] ),
    .Q(\alu_out_q[21] ));
 sky130_fd_sc_hd__dfxtp_2 _26437_ (.CLK(clk),
    .D(\alu_out[22] ),
    .Q(\alu_out_q[22] ));
 sky130_fd_sc_hd__dfxtp_2 _26438_ (.CLK(clk),
    .D(\alu_out[23] ),
    .Q(\alu_out_q[23] ));
 sky130_fd_sc_hd__dfxtp_2 _26439_ (.CLK(clk),
    .D(\alu_out[24] ),
    .Q(\alu_out_q[24] ));
 sky130_fd_sc_hd__dfxtp_2 _26440_ (.CLK(clk),
    .D(\alu_out[25] ),
    .Q(\alu_out_q[25] ));
 sky130_fd_sc_hd__dfxtp_2 _26441_ (.CLK(clk),
    .D(\alu_out[26] ),
    .Q(\alu_out_q[26] ));
 sky130_fd_sc_hd__dfxtp_2 _26442_ (.CLK(clk),
    .D(\alu_out[27] ),
    .Q(\alu_out_q[27] ));
 sky130_fd_sc_hd__dfxtp_2 _26443_ (.CLK(clk),
    .D(\alu_out[28] ),
    .Q(\alu_out_q[28] ));
 sky130_fd_sc_hd__dfxtp_2 _26444_ (.CLK(clk),
    .D(\alu_out[29] ),
    .Q(\alu_out_q[29] ));
 sky130_fd_sc_hd__dfxtp_2 _26445_ (.CLK(clk),
    .D(\alu_out[30] ),
    .Q(\alu_out_q[30] ));
 sky130_fd_sc_hd__dfxtp_2 _26446_ (.CLK(clk),
    .D(\alu_out[31] ),
    .Q(\alu_out_q[31] ));
 sky130_fd_sc_hd__dfxtp_2 _26447_ (.CLK(clk),
    .D(_00005_),
    .Q(is_lui_auipc_jal));
 sky130_fd_sc_hd__dfxtp_2 _26448_ (.CLK(clk),
    .D(_00006_),
    .Q(is_slti_blt_slt));
 sky130_fd_sc_hd__dfxtp_2 _26449_ (.CLK(clk),
    .D(_00007_),
    .Q(is_sltiu_bltu_sltu));
 sky130_fd_sc_hd__dfxtp_2 _26450_ (.CLK(clk),
    .D(_02591_),
    .Q(\alu_add_sub[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26451_ (.CLK(clk),
    .D(_02602_),
    .Q(\alu_add_sub[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26452_ (.CLK(clk),
    .D(_02613_),
    .Q(\alu_add_sub[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26453_ (.CLK(clk),
    .D(_02616_),
    .Q(\alu_add_sub[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26454_ (.CLK(clk),
    .D(_02617_),
    .Q(\alu_add_sub[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26455_ (.CLK(clk),
    .D(_02618_),
    .Q(\alu_add_sub[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26456_ (.CLK(clk),
    .D(_02619_),
    .Q(\alu_add_sub[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26457_ (.CLK(clk),
    .D(_02620_),
    .Q(\alu_add_sub[7] ));
 sky130_fd_sc_hd__dfxtp_2 _26458_ (.CLK(clk),
    .D(_02621_),
    .Q(\alu_add_sub[8] ));
 sky130_fd_sc_hd__dfxtp_2 _26459_ (.CLK(clk),
    .D(_02622_),
    .Q(\alu_add_sub[9] ));
 sky130_fd_sc_hd__dfxtp_2 _26460_ (.CLK(clk),
    .D(_02592_),
    .Q(\alu_add_sub[10] ));
 sky130_fd_sc_hd__dfxtp_2 _26461_ (.CLK(clk),
    .D(_02593_),
    .Q(\alu_add_sub[11] ));
 sky130_fd_sc_hd__dfxtp_2 _26462_ (.CLK(clk),
    .D(_02594_),
    .Q(\alu_add_sub[12] ));
 sky130_fd_sc_hd__dfxtp_2 _26463_ (.CLK(clk),
    .D(_02595_),
    .Q(\alu_add_sub[13] ));
 sky130_fd_sc_hd__dfxtp_2 _26464_ (.CLK(clk),
    .D(_02596_),
    .Q(\alu_add_sub[14] ));
 sky130_fd_sc_hd__dfxtp_2 _26465_ (.CLK(clk),
    .D(_02597_),
    .Q(\alu_add_sub[15] ));
 sky130_fd_sc_hd__dfxtp_2 _26466_ (.CLK(clk),
    .D(_02598_),
    .Q(\alu_add_sub[16] ));
 sky130_fd_sc_hd__dfxtp_2 _26467_ (.CLK(clk),
    .D(_02599_),
    .Q(\alu_add_sub[17] ));
 sky130_fd_sc_hd__dfxtp_2 _26468_ (.CLK(clk),
    .D(_02600_),
    .Q(\alu_add_sub[18] ));
 sky130_fd_sc_hd__dfxtp_2 _26469_ (.CLK(clk),
    .D(_02601_),
    .Q(\alu_add_sub[19] ));
 sky130_fd_sc_hd__dfxtp_2 _26470_ (.CLK(clk),
    .D(_02603_),
    .Q(\alu_add_sub[20] ));
 sky130_fd_sc_hd__dfxtp_2 _26471_ (.CLK(clk),
    .D(_02604_),
    .Q(\alu_add_sub[21] ));
 sky130_fd_sc_hd__dfxtp_2 _26472_ (.CLK(clk),
    .D(_02605_),
    .Q(\alu_add_sub[22] ));
 sky130_fd_sc_hd__dfxtp_2 _26473_ (.CLK(clk),
    .D(_02606_),
    .Q(\alu_add_sub[23] ));
 sky130_fd_sc_hd__dfxtp_2 _26474_ (.CLK(clk),
    .D(_02607_),
    .Q(\alu_add_sub[24] ));
 sky130_fd_sc_hd__dfxtp_2 _26475_ (.CLK(clk),
    .D(_02608_),
    .Q(\alu_add_sub[25] ));
 sky130_fd_sc_hd__dfxtp_2 _26476_ (.CLK(clk),
    .D(_02609_),
    .Q(\alu_add_sub[26] ));
 sky130_fd_sc_hd__dfxtp_2 _26477_ (.CLK(clk),
    .D(_02610_),
    .Q(\alu_add_sub[27] ));
 sky130_fd_sc_hd__dfxtp_2 _26478_ (.CLK(clk),
    .D(_02611_),
    .Q(\alu_add_sub[28] ));
 sky130_fd_sc_hd__dfxtp_2 _26479_ (.CLK(clk),
    .D(_02612_),
    .Q(\alu_add_sub[29] ));
 sky130_fd_sc_hd__dfxtp_2 _26480_ (.CLK(clk),
    .D(_02614_),
    .Q(\alu_add_sub[30] ));
 sky130_fd_sc_hd__dfxtp_2 _26481_ (.CLK(clk),
    .D(_02615_),
    .Q(\alu_add_sub[31] ));
 sky130_fd_sc_hd__dfxtp_2 _26482_ (.CLK(clk),
    .D(_12983_),
    .Q(\alu_shl[16] ));
 sky130_fd_sc_hd__dfxtp_2 _26483_ (.CLK(clk),
    .D(_12984_),
    .Q(\alu_shl[17] ));
 sky130_fd_sc_hd__dfxtp_2 _26484_ (.CLK(clk),
    .D(_12985_),
    .Q(\alu_shl[18] ));
 sky130_fd_sc_hd__dfxtp_2 _26485_ (.CLK(clk),
    .D(_12986_),
    .Q(\alu_shl[19] ));
 sky130_fd_sc_hd__dfxtp_2 _26486_ (.CLK(clk),
    .D(_12987_),
    .Q(\alu_shl[20] ));
 sky130_fd_sc_hd__dfxtp_2 _26487_ (.CLK(clk),
    .D(_12988_),
    .Q(\alu_shl[21] ));
 sky130_fd_sc_hd__dfxtp_2 _26488_ (.CLK(clk),
    .D(_12989_),
    .Q(\alu_shl[22] ));
 sky130_fd_sc_hd__dfxtp_2 _26489_ (.CLK(clk),
    .D(_12990_),
    .Q(\alu_shl[23] ));
 sky130_fd_sc_hd__dfxtp_2 _26490_ (.CLK(clk),
    .D(_12991_),
    .Q(\alu_shl[24] ));
 sky130_fd_sc_hd__dfxtp_2 _26491_ (.CLK(clk),
    .D(_12992_),
    .Q(\alu_shl[25] ));
 sky130_fd_sc_hd__dfxtp_2 _26492_ (.CLK(clk),
    .D(_12993_),
    .Q(\alu_shl[26] ));
 sky130_fd_sc_hd__dfxtp_2 _26493_ (.CLK(clk),
    .D(_12994_),
    .Q(\alu_shl[27] ));
 sky130_fd_sc_hd__dfxtp_2 _26494_ (.CLK(clk),
    .D(_12995_),
    .Q(\alu_shl[28] ));
 sky130_fd_sc_hd__dfxtp_2 _26495_ (.CLK(clk),
    .D(_12996_),
    .Q(\alu_shl[29] ));
 sky130_fd_sc_hd__dfxtp_2 _26496_ (.CLK(clk),
    .D(_12997_),
    .Q(\alu_shl[30] ));
 sky130_fd_sc_hd__dfxtp_2 _26497_ (.CLK(clk),
    .D(_12998_),
    .Q(\alu_shl[31] ));
 sky130_fd_sc_hd__dfxtp_2 _26498_ (.CLK(clk),
    .D(_12999_),
    .Q(\alu_shr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26499_ (.CLK(clk),
    .D(_13010_),
    .Q(\alu_shr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26500_ (.CLK(clk),
    .D(_13021_),
    .Q(\alu_shr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26501_ (.CLK(clk),
    .D(_13024_),
    .Q(\alu_shr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26502_ (.CLK(clk),
    .D(_13025_),
    .Q(\alu_shr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26503_ (.CLK(clk),
    .D(_13026_),
    .Q(\alu_shr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26504_ (.CLK(clk),
    .D(_13027_),
    .Q(\alu_shr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26505_ (.CLK(clk),
    .D(_13028_),
    .Q(\alu_shr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _26506_ (.CLK(clk),
    .D(_13029_),
    .Q(\alu_shr[8] ));
 sky130_fd_sc_hd__dfxtp_2 _26507_ (.CLK(clk),
    .D(_13030_),
    .Q(\alu_shr[9] ));
 sky130_fd_sc_hd__dfxtp_2 _26508_ (.CLK(clk),
    .D(_13000_),
    .Q(\alu_shr[10] ));
 sky130_fd_sc_hd__dfxtp_2 _26509_ (.CLK(clk),
    .D(_13001_),
    .Q(\alu_shr[11] ));
 sky130_fd_sc_hd__dfxtp_2 _26510_ (.CLK(clk),
    .D(_13002_),
    .Q(\alu_shr[12] ));
 sky130_fd_sc_hd__dfxtp_2 _26511_ (.CLK(clk),
    .D(_13003_),
    .Q(\alu_shr[13] ));
 sky130_fd_sc_hd__dfxtp_2 _26512_ (.CLK(clk),
    .D(_13004_),
    .Q(\alu_shr[14] ));
 sky130_fd_sc_hd__dfxtp_2 _26513_ (.CLK(clk),
    .D(_13005_),
    .Q(\alu_shr[15] ));
 sky130_fd_sc_hd__dfxtp_2 _26514_ (.CLK(clk),
    .D(_13006_),
    .Q(\alu_shr[16] ));
 sky130_fd_sc_hd__dfxtp_2 _26515_ (.CLK(clk),
    .D(_13007_),
    .Q(\alu_shr[17] ));
 sky130_fd_sc_hd__dfxtp_2 _26516_ (.CLK(clk),
    .D(_13008_),
    .Q(\alu_shr[18] ));
 sky130_fd_sc_hd__dfxtp_2 _26517_ (.CLK(clk),
    .D(_13009_),
    .Q(\alu_shr[19] ));
 sky130_fd_sc_hd__dfxtp_2 _26518_ (.CLK(clk),
    .D(_13011_),
    .Q(\alu_shr[20] ));
 sky130_fd_sc_hd__dfxtp_2 _26519_ (.CLK(clk),
    .D(_13012_),
    .Q(\alu_shr[21] ));
 sky130_fd_sc_hd__dfxtp_2 _26520_ (.CLK(clk),
    .D(_13013_),
    .Q(\alu_shr[22] ));
 sky130_fd_sc_hd__dfxtp_2 _26521_ (.CLK(clk),
    .D(_13014_),
    .Q(\alu_shr[23] ));
 sky130_fd_sc_hd__dfxtp_2 _26522_ (.CLK(clk),
    .D(_13015_),
    .Q(\alu_shr[24] ));
 sky130_fd_sc_hd__dfxtp_2 _26523_ (.CLK(clk),
    .D(_13016_),
    .Q(\alu_shr[25] ));
 sky130_fd_sc_hd__dfxtp_2 _26524_ (.CLK(clk),
    .D(_13017_),
    .Q(\alu_shr[26] ));
 sky130_fd_sc_hd__dfxtp_2 _26525_ (.CLK(clk),
    .D(_13018_),
    .Q(\alu_shr[27] ));
 sky130_fd_sc_hd__dfxtp_2 _26526_ (.CLK(clk),
    .D(_13019_),
    .Q(\alu_shr[28] ));
 sky130_fd_sc_hd__dfxtp_2 _26527_ (.CLK(clk),
    .D(_13020_),
    .Q(\alu_shr[29] ));
 sky130_fd_sc_hd__dfxtp_2 _26528_ (.CLK(clk),
    .D(_13022_),
    .Q(\alu_shr[30] ));
 sky130_fd_sc_hd__dfxtp_2 _26529_ (.CLK(clk),
    .D(_13023_),
    .Q(\alu_shr[31] ));
 sky130_fd_sc_hd__dfxtp_2 _26530_ (.CLK(clk),
    .D(_00000_),
    .Q(alu_eq));
 sky130_fd_sc_hd__dfxtp_2 _26531_ (.CLK(clk),
    .D(_00002_),
    .Q(alu_ltu));
 sky130_fd_sc_hd__dfxtp_2 _26532_ (.CLK(clk),
    .D(_00001_),
    .Q(alu_lts));
 sky130_fd_sc_hd__dfxtp_2 _26533_ (.CLK(clk),
    .D(_02623_),
    .Q(\pcpi_mul.rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26534_ (.CLK(clk),
    .D(_02624_),
    .Q(\pcpi_mul.rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26535_ (.CLK(clk),
    .D(_02625_),
    .Q(\pcpi_mul.rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26536_ (.CLK(clk),
    .D(_02626_),
    .Q(\pcpi_mul.rd[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26537_ (.CLK(clk),
    .D(_02627_),
    .Q(\pcpi_mul.rd[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26538_ (.CLK(clk),
    .D(_02628_),
    .Q(\pcpi_mul.rd[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26539_ (.CLK(clk),
    .D(_02683_),
    .Q(\pcpi_mul.rd[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26540_ (.CLK(clk),
    .D(_02684_),
    .Q(\pcpi_mul.rd[7] ));
 sky130_fd_sc_hd__dfxtp_2 _26541_ (.CLK(clk),
    .D(_02685_),
    .Q(\pcpi_mul.rd[8] ));
 sky130_fd_sc_hd__dfxtp_2 _26542_ (.CLK(clk),
    .D(_02686_),
    .Q(\pcpi_mul.rd[9] ));
 sky130_fd_sc_hd__dfxtp_2 _26543_ (.CLK(clk),
    .D(_02629_),
    .Q(\pcpi_mul.rd[10] ));
 sky130_fd_sc_hd__dfxtp_2 _26544_ (.CLK(clk),
    .D(_02630_),
    .Q(\pcpi_mul.rd[11] ));
 sky130_fd_sc_hd__dfxtp_2 _26545_ (.CLK(clk),
    .D(_02631_),
    .Q(\pcpi_mul.rd[12] ));
 sky130_fd_sc_hd__dfxtp_2 _26546_ (.CLK(clk),
    .D(_02632_),
    .Q(\pcpi_mul.rd[13] ));
 sky130_fd_sc_hd__dfxtp_2 _26547_ (.CLK(clk),
    .D(_02633_),
    .Q(\pcpi_mul.rd[14] ));
 sky130_fd_sc_hd__dfxtp_2 _26548_ (.CLK(clk),
    .D(_02634_),
    .Q(\pcpi_mul.rd[15] ));
 sky130_fd_sc_hd__dfxtp_2 _26549_ (.CLK(clk),
    .D(_02635_),
    .Q(\pcpi_mul.rd[16] ));
 sky130_fd_sc_hd__dfxtp_2 _26550_ (.CLK(clk),
    .D(_02636_),
    .Q(\pcpi_mul.rd[17] ));
 sky130_fd_sc_hd__dfxtp_2 _26551_ (.CLK(clk),
    .D(_02637_),
    .Q(\pcpi_mul.rd[18] ));
 sky130_fd_sc_hd__dfxtp_2 _26552_ (.CLK(clk),
    .D(_02638_),
    .Q(\pcpi_mul.rd[19] ));
 sky130_fd_sc_hd__dfxtp_2 _26553_ (.CLK(clk),
    .D(_02639_),
    .Q(\pcpi_mul.rd[20] ));
 sky130_fd_sc_hd__dfxtp_2 _26554_ (.CLK(clk),
    .D(_02640_),
    .Q(\pcpi_mul.rd[21] ));
 sky130_fd_sc_hd__dfxtp_2 _26555_ (.CLK(clk),
    .D(_02641_),
    .Q(\pcpi_mul.rd[22] ));
 sky130_fd_sc_hd__dfxtp_2 _26556_ (.CLK(clk),
    .D(_02642_),
    .Q(\pcpi_mul.rd[23] ));
 sky130_fd_sc_hd__dfxtp_2 _26557_ (.CLK(clk),
    .D(_02643_),
    .Q(\pcpi_mul.rd[24] ));
 sky130_fd_sc_hd__dfxtp_2 _26558_ (.CLK(clk),
    .D(_02644_),
    .Q(\pcpi_mul.rd[25] ));
 sky130_fd_sc_hd__dfxtp_2 _26559_ (.CLK(clk),
    .D(_02645_),
    .Q(\pcpi_mul.rd[26] ));
 sky130_fd_sc_hd__dfxtp_2 _26560_ (.CLK(clk),
    .D(_02646_),
    .Q(\pcpi_mul.rd[27] ));
 sky130_fd_sc_hd__dfxtp_2 _26561_ (.CLK(clk),
    .D(_02647_),
    .Q(\pcpi_mul.rd[28] ));
 sky130_fd_sc_hd__dfxtp_2 _26562_ (.CLK(clk),
    .D(_02648_),
    .Q(\pcpi_mul.rd[29] ));
 sky130_fd_sc_hd__dfxtp_2 _26563_ (.CLK(clk),
    .D(_02649_),
    .Q(\pcpi_mul.rd[30] ));
 sky130_fd_sc_hd__dfxtp_2 _26564_ (.CLK(clk),
    .D(_02650_),
    .Q(\pcpi_mul.rd[31] ));
 sky130_fd_sc_hd__dfxtp_2 _26565_ (.CLK(clk),
    .D(_02651_),
    .Q(\pcpi_mul.rd[32] ));
 sky130_fd_sc_hd__dfxtp_2 _26566_ (.CLK(clk),
    .D(_02652_),
    .Q(\pcpi_mul.rd[33] ));
 sky130_fd_sc_hd__dfxtp_2 _26567_ (.CLK(clk),
    .D(_02653_),
    .Q(\pcpi_mul.rd[34] ));
 sky130_fd_sc_hd__dfxtp_2 _26568_ (.CLK(clk),
    .D(_02654_),
    .Q(\pcpi_mul.rd[35] ));
 sky130_fd_sc_hd__dfxtp_2 _26569_ (.CLK(clk),
    .D(_02655_),
    .Q(\pcpi_mul.rd[36] ));
 sky130_fd_sc_hd__dfxtp_2 _26570_ (.CLK(clk),
    .D(_02656_),
    .Q(\pcpi_mul.rd[37] ));
 sky130_fd_sc_hd__dfxtp_2 _26571_ (.CLK(clk),
    .D(_02657_),
    .Q(\pcpi_mul.rd[38] ));
 sky130_fd_sc_hd__dfxtp_2 _26572_ (.CLK(clk),
    .D(_02658_),
    .Q(\pcpi_mul.rd[39] ));
 sky130_fd_sc_hd__dfxtp_2 _26573_ (.CLK(clk),
    .D(_02659_),
    .Q(\pcpi_mul.rd[40] ));
 sky130_fd_sc_hd__dfxtp_2 _26574_ (.CLK(clk),
    .D(_02660_),
    .Q(\pcpi_mul.rd[41] ));
 sky130_fd_sc_hd__dfxtp_2 _26575_ (.CLK(clk),
    .D(_02661_),
    .Q(\pcpi_mul.rd[42] ));
 sky130_fd_sc_hd__dfxtp_2 _26576_ (.CLK(clk),
    .D(_02662_),
    .Q(\pcpi_mul.rd[43] ));
 sky130_fd_sc_hd__dfxtp_2 _26577_ (.CLK(clk),
    .D(_02663_),
    .Q(\pcpi_mul.rd[44] ));
 sky130_fd_sc_hd__dfxtp_2 _26578_ (.CLK(clk),
    .D(_02664_),
    .Q(\pcpi_mul.rd[45] ));
 sky130_fd_sc_hd__dfxtp_2 _26579_ (.CLK(clk),
    .D(_02665_),
    .Q(\pcpi_mul.rd[46] ));
 sky130_fd_sc_hd__dfxtp_2 _26580_ (.CLK(clk),
    .D(_02666_),
    .Q(\pcpi_mul.rd[47] ));
 sky130_fd_sc_hd__dfxtp_2 _26581_ (.CLK(clk),
    .D(_02667_),
    .Q(\pcpi_mul.rd[48] ));
 sky130_fd_sc_hd__dfxtp_2 _26582_ (.CLK(clk),
    .D(_02668_),
    .Q(\pcpi_mul.rd[49] ));
 sky130_fd_sc_hd__dfxtp_2 _26583_ (.CLK(clk),
    .D(_02669_),
    .Q(\pcpi_mul.rd[50] ));
 sky130_fd_sc_hd__dfxtp_2 _26584_ (.CLK(clk),
    .D(_02670_),
    .Q(\pcpi_mul.rd[51] ));
 sky130_fd_sc_hd__dfxtp_2 _26585_ (.CLK(clk),
    .D(_02671_),
    .Q(\pcpi_mul.rd[52] ));
 sky130_fd_sc_hd__dfxtp_2 _26586_ (.CLK(clk),
    .D(_02672_),
    .Q(\pcpi_mul.rd[53] ));
 sky130_fd_sc_hd__dfxtp_2 _26587_ (.CLK(clk),
    .D(_02673_),
    .Q(\pcpi_mul.rd[54] ));
 sky130_fd_sc_hd__dfxtp_2 _26588_ (.CLK(clk),
    .D(_02674_),
    .Q(\pcpi_mul.rd[55] ));
 sky130_fd_sc_hd__dfxtp_2 _26589_ (.CLK(clk),
    .D(_02675_),
    .Q(\pcpi_mul.rd[56] ));
 sky130_fd_sc_hd__dfxtp_2 _26590_ (.CLK(clk),
    .D(_02676_),
    .Q(\pcpi_mul.rd[57] ));
 sky130_fd_sc_hd__dfxtp_2 _26591_ (.CLK(clk),
    .D(_02677_),
    .Q(\pcpi_mul.rd[58] ));
 sky130_fd_sc_hd__dfxtp_2 _26592_ (.CLK(clk),
    .D(_02678_),
    .Q(\pcpi_mul.rd[59] ));
 sky130_fd_sc_hd__dfxtp_2 _26593_ (.CLK(clk),
    .D(_02679_),
    .Q(\pcpi_mul.rd[60] ));
 sky130_fd_sc_hd__dfxtp_2 _26594_ (.CLK(clk),
    .D(_02680_),
    .Q(\pcpi_mul.rd[61] ));
 sky130_fd_sc_hd__dfxtp_2 _26595_ (.CLK(clk),
    .D(_02681_),
    .Q(\pcpi_mul.rd[62] ));
 sky130_fd_sc_hd__dfxtp_2 _26596_ (.CLK(clk),
    .D(_02682_),
    .Q(\pcpi_mul.rd[63] ));
 sky130_fd_sc_hd__dfxtp_2 _26597_ (.CLK(clk),
    .D(\pcpi_mul.instr_any_mulh ),
    .Q(\pcpi_mul.shift_out ));
 sky130_fd_sc_hd__dfxtp_2 _26598_ (.CLK(clk),
    .D(_00038_),
    .Q(\cpu_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26599_ (.CLK(clk),
    .D(_00039_),
    .Q(\cpu_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26600_ (.CLK(clk),
    .D(_00040_),
    .Q(\cpu_state[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26601_ (.CLK(clk),
    .D(_00041_),
    .Q(\cpu_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26602_ (.CLK(clk),
    .D(_00042_),
    .Q(\cpu_state[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26603_ (.CLK(clk),
    .D(_00043_),
    .Q(\cpu_state[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26604_ (.CLK(clk),
    .D(_00044_),
    .Q(\cpu_state[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26605_ (.CLK(clk),
    .D(_02771_),
    .Q(\cpuregs[8][0] ));
 sky130_fd_sc_hd__dfxtp_2 _26606_ (.CLK(clk),
    .D(_02772_),
    .Q(\cpuregs[8][1] ));
 sky130_fd_sc_hd__dfxtp_2 _26607_ (.CLK(clk),
    .D(_02773_),
    .Q(\cpuregs[8][2] ));
 sky130_fd_sc_hd__dfxtp_2 _26608_ (.CLK(clk),
    .D(_02774_),
    .Q(\cpuregs[8][3] ));
 sky130_fd_sc_hd__dfxtp_2 _26609_ (.CLK(clk),
    .D(_02775_),
    .Q(\cpuregs[8][4] ));
 sky130_fd_sc_hd__dfxtp_2 _26610_ (.CLK(clk),
    .D(_02776_),
    .Q(\cpuregs[8][5] ));
 sky130_fd_sc_hd__dfxtp_2 _26611_ (.CLK(clk),
    .D(_02777_),
    .Q(\cpuregs[8][6] ));
 sky130_fd_sc_hd__dfxtp_2 _26612_ (.CLK(clk),
    .D(_02778_),
    .Q(\cpuregs[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _26613_ (.CLK(clk),
    .D(_02779_),
    .Q(\cpuregs[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _26614_ (.CLK(clk),
    .D(_02780_),
    .Q(\cpuregs[8][9] ));
 sky130_fd_sc_hd__dfxtp_2 _26615_ (.CLK(clk),
    .D(_02781_),
    .Q(\cpuregs[8][10] ));
 sky130_fd_sc_hd__dfxtp_2 _26616_ (.CLK(clk),
    .D(_02782_),
    .Q(\cpuregs[8][11] ));
 sky130_fd_sc_hd__dfxtp_2 _26617_ (.CLK(clk),
    .D(_02783_),
    .Q(\cpuregs[8][12] ));
 sky130_fd_sc_hd__dfxtp_2 _26618_ (.CLK(clk),
    .D(_02784_),
    .Q(\cpuregs[8][13] ));
 sky130_fd_sc_hd__dfxtp_2 _26619_ (.CLK(clk),
    .D(_02785_),
    .Q(\cpuregs[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _26620_ (.CLK(clk),
    .D(_02786_),
    .Q(\cpuregs[8][15] ));
 sky130_fd_sc_hd__dfxtp_2 _26621_ (.CLK(clk),
    .D(_02787_),
    .Q(\cpuregs[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _26622_ (.CLK(clk),
    .D(_02788_),
    .Q(\cpuregs[8][17] ));
 sky130_fd_sc_hd__dfxtp_2 _26623_ (.CLK(clk),
    .D(_02789_),
    .Q(\cpuregs[8][18] ));
 sky130_fd_sc_hd__dfxtp_2 _26624_ (.CLK(clk),
    .D(_02790_),
    .Q(\cpuregs[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _26625_ (.CLK(clk),
    .D(_02791_),
    .Q(\cpuregs[8][20] ));
 sky130_fd_sc_hd__dfxtp_2 _26626_ (.CLK(clk),
    .D(_02792_),
    .Q(\cpuregs[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _26627_ (.CLK(clk),
    .D(_02793_),
    .Q(\cpuregs[8][22] ));
 sky130_fd_sc_hd__dfxtp_2 _26628_ (.CLK(clk),
    .D(_02794_),
    .Q(\cpuregs[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _26629_ (.CLK(clk),
    .D(_02795_),
    .Q(\cpuregs[8][24] ));
 sky130_fd_sc_hd__dfxtp_2 _26630_ (.CLK(clk),
    .D(_02796_),
    .Q(\cpuregs[8][25] ));
 sky130_fd_sc_hd__dfxtp_2 _26631_ (.CLK(clk),
    .D(_02797_),
    .Q(\cpuregs[8][26] ));
 sky130_fd_sc_hd__dfxtp_2 _26632_ (.CLK(clk),
    .D(_02798_),
    .Q(\cpuregs[8][27] ));
 sky130_fd_sc_hd__dfxtp_2 _26633_ (.CLK(clk),
    .D(_02799_),
    .Q(\cpuregs[8][28] ));
 sky130_fd_sc_hd__dfxtp_2 _26634_ (.CLK(clk),
    .D(_02800_),
    .Q(\cpuregs[8][29] ));
 sky130_fd_sc_hd__dfxtp_2 _26635_ (.CLK(clk),
    .D(_02801_),
    .Q(\cpuregs[8][30] ));
 sky130_fd_sc_hd__dfxtp_2 _26636_ (.CLK(clk),
    .D(_02802_),
    .Q(\cpuregs[8][31] ));
 sky130_fd_sc_hd__dfxtp_2 _26637_ (.CLK(clk),
    .D(_02803_),
    .Q(\cpuregs[14][0] ));
 sky130_fd_sc_hd__dfxtp_2 _26638_ (.CLK(clk),
    .D(_02804_),
    .Q(\cpuregs[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _26639_ (.CLK(clk),
    .D(_02805_),
    .Q(\cpuregs[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _26640_ (.CLK(clk),
    .D(_02806_),
    .Q(\cpuregs[14][3] ));
 sky130_fd_sc_hd__dfxtp_2 _26641_ (.CLK(clk),
    .D(_02807_),
    .Q(\cpuregs[14][4] ));
 sky130_fd_sc_hd__dfxtp_2 _26642_ (.CLK(clk),
    .D(_02808_),
    .Q(\cpuregs[14][5] ));
 sky130_fd_sc_hd__dfxtp_2 _26643_ (.CLK(clk),
    .D(_02809_),
    .Q(\cpuregs[14][6] ));
 sky130_fd_sc_hd__dfxtp_2 _26644_ (.CLK(clk),
    .D(_02810_),
    .Q(\cpuregs[14][7] ));
 sky130_fd_sc_hd__dfxtp_2 _26645_ (.CLK(clk),
    .D(_02811_),
    .Q(\cpuregs[14][8] ));
 sky130_fd_sc_hd__dfxtp_2 _26646_ (.CLK(clk),
    .D(_02812_),
    .Q(\cpuregs[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _26647_ (.CLK(clk),
    .D(_02813_),
    .Q(\cpuregs[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _26648_ (.CLK(clk),
    .D(_02814_),
    .Q(\cpuregs[14][11] ));
 sky130_fd_sc_hd__dfxtp_2 _26649_ (.CLK(clk),
    .D(_02815_),
    .Q(\cpuregs[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _26650_ (.CLK(clk),
    .D(_02816_),
    .Q(\cpuregs[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _26651_ (.CLK(clk),
    .D(_02817_),
    .Q(\cpuregs[14][14] ));
 sky130_fd_sc_hd__dfxtp_2 _26652_ (.CLK(clk),
    .D(_02818_),
    .Q(\cpuregs[14][15] ));
 sky130_fd_sc_hd__dfxtp_2 _26653_ (.CLK(clk),
    .D(_02819_),
    .Q(\cpuregs[14][16] ));
 sky130_fd_sc_hd__dfxtp_2 _26654_ (.CLK(clk),
    .D(_02820_),
    .Q(\cpuregs[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _26655_ (.CLK(clk),
    .D(_02821_),
    .Q(\cpuregs[14][18] ));
 sky130_fd_sc_hd__dfxtp_2 _26656_ (.CLK(clk),
    .D(_02822_),
    .Q(\cpuregs[14][19] ));
 sky130_fd_sc_hd__dfxtp_2 _26657_ (.CLK(clk),
    .D(_02823_),
    .Q(\cpuregs[14][20] ));
 sky130_fd_sc_hd__dfxtp_2 _26658_ (.CLK(clk),
    .D(_02824_),
    .Q(\cpuregs[14][21] ));
 sky130_fd_sc_hd__dfxtp_2 _26659_ (.CLK(clk),
    .D(_02825_),
    .Q(\cpuregs[14][22] ));
 sky130_fd_sc_hd__dfxtp_2 _26660_ (.CLK(clk),
    .D(_02826_),
    .Q(\cpuregs[14][23] ));
 sky130_fd_sc_hd__dfxtp_2 _26661_ (.CLK(clk),
    .D(_02827_),
    .Q(\cpuregs[14][24] ));
 sky130_fd_sc_hd__dfxtp_2 _26662_ (.CLK(clk),
    .D(_02828_),
    .Q(\cpuregs[14][25] ));
 sky130_fd_sc_hd__dfxtp_2 _26663_ (.CLK(clk),
    .D(_02829_),
    .Q(\cpuregs[14][26] ));
 sky130_fd_sc_hd__dfxtp_2 _26664_ (.CLK(clk),
    .D(_02830_),
    .Q(\cpuregs[14][27] ));
 sky130_fd_sc_hd__dfxtp_2 _26665_ (.CLK(clk),
    .D(_02831_),
    .Q(\cpuregs[14][28] ));
 sky130_fd_sc_hd__dfxtp_2 _26666_ (.CLK(clk),
    .D(_02832_),
    .Q(\cpuregs[14][29] ));
 sky130_fd_sc_hd__dfxtp_2 _26667_ (.CLK(clk),
    .D(_02833_),
    .Q(\cpuregs[14][30] ));
 sky130_fd_sc_hd__dfxtp_2 _26668_ (.CLK(clk),
    .D(_02834_),
    .Q(\cpuregs[14][31] ));
 sky130_fd_sc_hd__dfxtp_2 _26669_ (.CLK(clk),
    .D(_02835_),
    .Q(\cpuregs[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _26670_ (.CLK(clk),
    .D(_02836_),
    .Q(\cpuregs[0][1] ));
 sky130_fd_sc_hd__dfxtp_2 _26671_ (.CLK(clk),
    .D(_02837_),
    .Q(\cpuregs[0][2] ));
 sky130_fd_sc_hd__dfxtp_2 _26672_ (.CLK(clk),
    .D(_02838_),
    .Q(\cpuregs[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _26673_ (.CLK(clk),
    .D(_02839_),
    .Q(\cpuregs[0][4] ));
 sky130_fd_sc_hd__dfxtp_2 _26674_ (.CLK(clk),
    .D(_02840_),
    .Q(\cpuregs[0][5] ));
 sky130_fd_sc_hd__dfxtp_2 _26675_ (.CLK(clk),
    .D(_02841_),
    .Q(\cpuregs[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _26676_ (.CLK(clk),
    .D(_02842_),
    .Q(\cpuregs[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _26677_ (.CLK(clk),
    .D(_02843_),
    .Q(\cpuregs[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _26678_ (.CLK(clk),
    .D(_02844_),
    .Q(\cpuregs[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _26679_ (.CLK(clk),
    .D(_02845_),
    .Q(\cpuregs[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _26680_ (.CLK(clk),
    .D(_02846_),
    .Q(\cpuregs[0][11] ));
 sky130_fd_sc_hd__dfxtp_2 _26681_ (.CLK(clk),
    .D(_02847_),
    .Q(\cpuregs[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _26682_ (.CLK(clk),
    .D(_02848_),
    .Q(\cpuregs[0][13] ));
 sky130_fd_sc_hd__dfxtp_2 _26683_ (.CLK(clk),
    .D(_02849_),
    .Q(\cpuregs[0][14] ));
 sky130_fd_sc_hd__dfxtp_2 _26684_ (.CLK(clk),
    .D(_02850_),
    .Q(\cpuregs[0][15] ));
 sky130_fd_sc_hd__dfxtp_2 _26685_ (.CLK(clk),
    .D(_02851_),
    .Q(\cpuregs[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _26686_ (.CLK(clk),
    .D(_02852_),
    .Q(\cpuregs[0][17] ));
 sky130_fd_sc_hd__dfxtp_2 _26687_ (.CLK(clk),
    .D(_02853_),
    .Q(\cpuregs[0][18] ));
 sky130_fd_sc_hd__dfxtp_2 _26688_ (.CLK(clk),
    .D(_02854_),
    .Q(\cpuregs[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _26689_ (.CLK(clk),
    .D(_02855_),
    .Q(\cpuregs[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _26690_ (.CLK(clk),
    .D(_02856_),
    .Q(\cpuregs[0][21] ));
 sky130_fd_sc_hd__dfxtp_2 _26691_ (.CLK(clk),
    .D(_02857_),
    .Q(\cpuregs[0][22] ));
 sky130_fd_sc_hd__dfxtp_2 _26692_ (.CLK(clk),
    .D(_02858_),
    .Q(\cpuregs[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _26693_ (.CLK(clk),
    .D(_02859_),
    .Q(\cpuregs[0][24] ));
 sky130_fd_sc_hd__dfxtp_2 _26694_ (.CLK(clk),
    .D(_02860_),
    .Q(\cpuregs[0][25] ));
 sky130_fd_sc_hd__dfxtp_2 _26695_ (.CLK(clk),
    .D(_02861_),
    .Q(\cpuregs[0][26] ));
 sky130_fd_sc_hd__dfxtp_2 _26696_ (.CLK(clk),
    .D(_02862_),
    .Q(\cpuregs[0][27] ));
 sky130_fd_sc_hd__dfxtp_2 _26697_ (.CLK(clk),
    .D(_02863_),
    .Q(\cpuregs[0][28] ));
 sky130_fd_sc_hd__dfxtp_2 _26698_ (.CLK(clk),
    .D(_02864_),
    .Q(\cpuregs[0][29] ));
 sky130_fd_sc_hd__dfxtp_2 _26699_ (.CLK(clk),
    .D(_02865_),
    .Q(\cpuregs[0][30] ));
 sky130_fd_sc_hd__dfxtp_2 _26700_ (.CLK(clk),
    .D(_02866_),
    .Q(\cpuregs[0][31] ));
 sky130_fd_sc_hd__dfxtp_2 _26701_ (.CLK(clk),
    .D(_02867_),
    .Q(\cpuregs[10][0] ));
 sky130_fd_sc_hd__dfxtp_2 _26702_ (.CLK(clk),
    .D(_02868_),
    .Q(\cpuregs[10][1] ));
 sky130_fd_sc_hd__dfxtp_2 _26703_ (.CLK(clk),
    .D(_02869_),
    .Q(\cpuregs[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _26704_ (.CLK(clk),
    .D(_02870_),
    .Q(\cpuregs[10][3] ));
 sky130_fd_sc_hd__dfxtp_2 _26705_ (.CLK(clk),
    .D(_02871_),
    .Q(\cpuregs[10][4] ));
 sky130_fd_sc_hd__dfxtp_2 _26706_ (.CLK(clk),
    .D(_02872_),
    .Q(\cpuregs[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _26707_ (.CLK(clk),
    .D(_02873_),
    .Q(\cpuregs[10][6] ));
 sky130_fd_sc_hd__dfxtp_2 _26708_ (.CLK(clk),
    .D(_02874_),
    .Q(\cpuregs[10][7] ));
 sky130_fd_sc_hd__dfxtp_2 _26709_ (.CLK(clk),
    .D(_02875_),
    .Q(\cpuregs[10][8] ));
 sky130_fd_sc_hd__dfxtp_2 _26710_ (.CLK(clk),
    .D(_02876_),
    .Q(\cpuregs[10][9] ));
 sky130_fd_sc_hd__dfxtp_2 _26711_ (.CLK(clk),
    .D(_02877_),
    .Q(\cpuregs[10][10] ));
 sky130_fd_sc_hd__dfxtp_2 _26712_ (.CLK(clk),
    .D(_02878_),
    .Q(\cpuregs[10][11] ));
 sky130_fd_sc_hd__dfxtp_2 _26713_ (.CLK(clk),
    .D(_02879_),
    .Q(\cpuregs[10][12] ));
 sky130_fd_sc_hd__dfxtp_2 _26714_ (.CLK(clk),
    .D(_02880_),
    .Q(\cpuregs[10][13] ));
 sky130_fd_sc_hd__dfxtp_2 _26715_ (.CLK(clk),
    .D(_02881_),
    .Q(\cpuregs[10][14] ));
 sky130_fd_sc_hd__dfxtp_2 _26716_ (.CLK(clk),
    .D(_02882_),
    .Q(\cpuregs[10][15] ));
 sky130_fd_sc_hd__dfxtp_2 _26717_ (.CLK(clk),
    .D(_02883_),
    .Q(\cpuregs[10][16] ));
 sky130_fd_sc_hd__dfxtp_2 _26718_ (.CLK(clk),
    .D(_02884_),
    .Q(\cpuregs[10][17] ));
 sky130_fd_sc_hd__dfxtp_2 _26719_ (.CLK(clk),
    .D(_02885_),
    .Q(\cpuregs[10][18] ));
 sky130_fd_sc_hd__dfxtp_2 _26720_ (.CLK(clk),
    .D(_02886_),
    .Q(\cpuregs[10][19] ));
 sky130_fd_sc_hd__dfxtp_2 _26721_ (.CLK(clk),
    .D(_02887_),
    .Q(\cpuregs[10][20] ));
 sky130_fd_sc_hd__dfxtp_2 _26722_ (.CLK(clk),
    .D(_02888_),
    .Q(\cpuregs[10][21] ));
 sky130_fd_sc_hd__dfxtp_2 _26723_ (.CLK(clk),
    .D(_02889_),
    .Q(\cpuregs[10][22] ));
 sky130_fd_sc_hd__dfxtp_2 _26724_ (.CLK(clk),
    .D(_02890_),
    .Q(\cpuregs[10][23] ));
 sky130_fd_sc_hd__dfxtp_2 _26725_ (.CLK(clk),
    .D(_02891_),
    .Q(\cpuregs[10][24] ));
 sky130_fd_sc_hd__dfxtp_2 _26726_ (.CLK(clk),
    .D(_02892_),
    .Q(\cpuregs[10][25] ));
 sky130_fd_sc_hd__dfxtp_2 _26727_ (.CLK(clk),
    .D(_02893_),
    .Q(\cpuregs[10][26] ));
 sky130_fd_sc_hd__dfxtp_2 _26728_ (.CLK(clk),
    .D(_02894_),
    .Q(\cpuregs[10][27] ));
 sky130_fd_sc_hd__dfxtp_2 _26729_ (.CLK(clk),
    .D(_02895_),
    .Q(\cpuregs[10][28] ));
 sky130_fd_sc_hd__dfxtp_2 _26730_ (.CLK(clk),
    .D(_02896_),
    .Q(\cpuregs[10][29] ));
 sky130_fd_sc_hd__dfxtp_2 _26731_ (.CLK(clk),
    .D(_02897_),
    .Q(\cpuregs[10][30] ));
 sky130_fd_sc_hd__dfxtp_2 _26732_ (.CLK(clk),
    .D(_02898_),
    .Q(\cpuregs[10][31] ));
 sky130_fd_sc_hd__dfxtp_2 _26733_ (.CLK(clk),
    .D(_02899_),
    .Q(\cpuregs[18][0] ));
 sky130_fd_sc_hd__dfxtp_2 _26734_ (.CLK(clk),
    .D(_02900_),
    .Q(\cpuregs[18][1] ));
 sky130_fd_sc_hd__dfxtp_2 _26735_ (.CLK(clk),
    .D(_02901_),
    .Q(\cpuregs[18][2] ));
 sky130_fd_sc_hd__dfxtp_2 _26736_ (.CLK(clk),
    .D(_02902_),
    .Q(\cpuregs[18][3] ));
 sky130_fd_sc_hd__dfxtp_2 _26737_ (.CLK(clk),
    .D(_02903_),
    .Q(\cpuregs[18][4] ));
 sky130_fd_sc_hd__dfxtp_2 _26738_ (.CLK(clk),
    .D(_02904_),
    .Q(\cpuregs[18][5] ));
 sky130_fd_sc_hd__dfxtp_2 _26739_ (.CLK(clk),
    .D(_02905_),
    .Q(\cpuregs[18][6] ));
 sky130_fd_sc_hd__dfxtp_2 _26740_ (.CLK(clk),
    .D(_02906_),
    .Q(\cpuregs[18][7] ));
 sky130_fd_sc_hd__dfxtp_2 _26741_ (.CLK(clk),
    .D(_02907_),
    .Q(\cpuregs[18][8] ));
 sky130_fd_sc_hd__dfxtp_2 _26742_ (.CLK(clk),
    .D(_02908_),
    .Q(\cpuregs[18][9] ));
 sky130_fd_sc_hd__dfxtp_2 _26743_ (.CLK(clk),
    .D(_02909_),
    .Q(\cpuregs[18][10] ));
 sky130_fd_sc_hd__dfxtp_2 _26744_ (.CLK(clk),
    .D(_02910_),
    .Q(\cpuregs[18][11] ));
 sky130_fd_sc_hd__dfxtp_2 _26745_ (.CLK(clk),
    .D(_02911_),
    .Q(\cpuregs[18][12] ));
 sky130_fd_sc_hd__dfxtp_2 _26746_ (.CLK(clk),
    .D(_02912_),
    .Q(\cpuregs[18][13] ));
 sky130_fd_sc_hd__dfxtp_2 _26747_ (.CLK(clk),
    .D(_02913_),
    .Q(\cpuregs[18][14] ));
 sky130_fd_sc_hd__dfxtp_2 _26748_ (.CLK(clk),
    .D(_02914_),
    .Q(\cpuregs[18][15] ));
 sky130_fd_sc_hd__dfxtp_2 _26749_ (.CLK(clk),
    .D(_02915_),
    .Q(\cpuregs[18][16] ));
 sky130_fd_sc_hd__dfxtp_2 _26750_ (.CLK(clk),
    .D(_02916_),
    .Q(\cpuregs[18][17] ));
 sky130_fd_sc_hd__dfxtp_2 _26751_ (.CLK(clk),
    .D(_02917_),
    .Q(\cpuregs[18][18] ));
 sky130_fd_sc_hd__dfxtp_2 _26752_ (.CLK(clk),
    .D(_02918_),
    .Q(\cpuregs[18][19] ));
 sky130_fd_sc_hd__dfxtp_2 _26753_ (.CLK(clk),
    .D(_02919_),
    .Q(\cpuregs[18][20] ));
 sky130_fd_sc_hd__dfxtp_2 _26754_ (.CLK(clk),
    .D(_02920_),
    .Q(\cpuregs[18][21] ));
 sky130_fd_sc_hd__dfxtp_2 _26755_ (.CLK(clk),
    .D(_02921_),
    .Q(\cpuregs[18][22] ));
 sky130_fd_sc_hd__dfxtp_2 _26756_ (.CLK(clk),
    .D(_02922_),
    .Q(\cpuregs[18][23] ));
 sky130_fd_sc_hd__dfxtp_2 _26757_ (.CLK(clk),
    .D(_02923_),
    .Q(\cpuregs[18][24] ));
 sky130_fd_sc_hd__dfxtp_2 _26758_ (.CLK(clk),
    .D(_02924_),
    .Q(\cpuregs[18][25] ));
 sky130_fd_sc_hd__dfxtp_2 _26759_ (.CLK(clk),
    .D(_02925_),
    .Q(\cpuregs[18][26] ));
 sky130_fd_sc_hd__dfxtp_2 _26760_ (.CLK(clk),
    .D(_02926_),
    .Q(\cpuregs[18][27] ));
 sky130_fd_sc_hd__dfxtp_2 _26761_ (.CLK(clk),
    .D(_02927_),
    .Q(\cpuregs[18][28] ));
 sky130_fd_sc_hd__dfxtp_2 _26762_ (.CLK(clk),
    .D(_02928_),
    .Q(\cpuregs[18][29] ));
 sky130_fd_sc_hd__dfxtp_2 _26763_ (.CLK(clk),
    .D(_02929_),
    .Q(\cpuregs[18][30] ));
 sky130_fd_sc_hd__dfxtp_2 _26764_ (.CLK(clk),
    .D(_02930_),
    .Q(\cpuregs[18][31] ));
 sky130_fd_sc_hd__dfxtp_2 _26765_ (.CLK(clk),
    .D(_02931_),
    .Q(\mem_rdata_q[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26766_ (.CLK(clk),
    .D(_02932_),
    .Q(\mem_rdata_q[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26767_ (.CLK(clk),
    .D(_02933_),
    .Q(\mem_rdata_q[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26768_ (.CLK(clk),
    .D(_02934_),
    .Q(\mem_rdata_q[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26769_ (.CLK(clk),
    .D(_02935_),
    .Q(\mem_rdata_q[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26770_ (.CLK(clk),
    .D(_02936_),
    .Q(\mem_rdata_q[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26771_ (.CLK(clk),
    .D(_02937_),
    .Q(\mem_rdata_q[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26772_ (.CLK(clk),
    .D(_02938_),
    .Q(\mem_rdata_q[7] ));
 sky130_fd_sc_hd__dfxtp_2 _26773_ (.CLK(clk),
    .D(_02939_),
    .Q(\mem_rdata_q[8] ));
 sky130_fd_sc_hd__dfxtp_2 _26774_ (.CLK(clk),
    .D(_02940_),
    .Q(\mem_rdata_q[9] ));
 sky130_fd_sc_hd__dfxtp_2 _26775_ (.CLK(clk),
    .D(_02941_),
    .Q(\mem_rdata_q[10] ));
 sky130_fd_sc_hd__dfxtp_2 _26776_ (.CLK(clk),
    .D(_02942_),
    .Q(\mem_rdata_q[11] ));
 sky130_fd_sc_hd__dfxtp_2 _26777_ (.CLK(clk),
    .D(_02943_),
    .Q(\mem_rdata_q[12] ));
 sky130_fd_sc_hd__dfxtp_2 _26778_ (.CLK(clk),
    .D(_02944_),
    .Q(\mem_rdata_q[13] ));
 sky130_fd_sc_hd__dfxtp_2 _26779_ (.CLK(clk),
    .D(_02945_),
    .Q(\mem_rdata_q[14] ));
 sky130_fd_sc_hd__dfxtp_2 _26780_ (.CLK(clk),
    .D(_02946_),
    .Q(\mem_rdata_q[15] ));
 sky130_fd_sc_hd__dfxtp_2 _26781_ (.CLK(clk),
    .D(_02947_),
    .Q(\mem_rdata_q[16] ));
 sky130_fd_sc_hd__dfxtp_2 _26782_ (.CLK(clk),
    .D(_02948_),
    .Q(\mem_rdata_q[17] ));
 sky130_fd_sc_hd__dfxtp_2 _26783_ (.CLK(clk),
    .D(_02949_),
    .Q(\mem_rdata_q[18] ));
 sky130_fd_sc_hd__dfxtp_2 _26784_ (.CLK(clk),
    .D(_02950_),
    .Q(\mem_rdata_q[19] ));
 sky130_fd_sc_hd__dfxtp_2 _26785_ (.CLK(clk),
    .D(_02951_),
    .Q(\mem_rdata_q[20] ));
 sky130_fd_sc_hd__dfxtp_2 _26786_ (.CLK(clk),
    .D(_02952_),
    .Q(\mem_rdata_q[21] ));
 sky130_fd_sc_hd__dfxtp_2 _26787_ (.CLK(clk),
    .D(_02953_),
    .Q(\mem_rdata_q[22] ));
 sky130_fd_sc_hd__dfxtp_2 _26788_ (.CLK(clk),
    .D(_02954_),
    .Q(\mem_rdata_q[23] ));
 sky130_fd_sc_hd__dfxtp_2 _26789_ (.CLK(clk),
    .D(_02955_),
    .Q(\mem_rdata_q[24] ));
 sky130_fd_sc_hd__dfxtp_2 _26790_ (.CLK(clk),
    .D(_02956_),
    .Q(\mem_rdata_q[25] ));
 sky130_fd_sc_hd__dfxtp_2 _26791_ (.CLK(clk),
    .D(_02957_),
    .Q(\mem_rdata_q[26] ));
 sky130_fd_sc_hd__dfxtp_2 _26792_ (.CLK(clk),
    .D(_02958_),
    .Q(\mem_rdata_q[27] ));
 sky130_fd_sc_hd__dfxtp_2 _26793_ (.CLK(clk),
    .D(_02959_),
    .Q(\mem_rdata_q[28] ));
 sky130_fd_sc_hd__dfxtp_2 _26794_ (.CLK(clk),
    .D(_02960_),
    .Q(\mem_rdata_q[29] ));
 sky130_fd_sc_hd__dfxtp_2 _26795_ (.CLK(clk),
    .D(_02961_),
    .Q(\mem_rdata_q[30] ));
 sky130_fd_sc_hd__dfxtp_2 _26796_ (.CLK(clk),
    .D(_02962_),
    .Q(\mem_rdata_q[31] ));
 sky130_fd_sc_hd__dfxtp_2 _26797_ (.CLK(clk),
    .D(_02963_),
    .Q(\cpuregs[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _26798_ (.CLK(clk),
    .D(_02964_),
    .Q(\cpuregs[2][1] ));
 sky130_fd_sc_hd__dfxtp_2 _26799_ (.CLK(clk),
    .D(_02965_),
    .Q(\cpuregs[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _26800_ (.CLK(clk),
    .D(_02966_),
    .Q(\cpuregs[2][3] ));
 sky130_fd_sc_hd__dfxtp_2 _26801_ (.CLK(clk),
    .D(_02967_),
    .Q(\cpuregs[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _26802_ (.CLK(clk),
    .D(_02968_),
    .Q(\cpuregs[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _26803_ (.CLK(clk),
    .D(_02969_),
    .Q(\cpuregs[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _26804_ (.CLK(clk),
    .D(_02970_),
    .Q(\cpuregs[2][7] ));
 sky130_fd_sc_hd__dfxtp_2 _26805_ (.CLK(clk),
    .D(_02971_),
    .Q(\cpuregs[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _26806_ (.CLK(clk),
    .D(_02972_),
    .Q(\cpuregs[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _26807_ (.CLK(clk),
    .D(_02973_),
    .Q(\cpuregs[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _26808_ (.CLK(clk),
    .D(_02974_),
    .Q(\cpuregs[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _26809_ (.CLK(clk),
    .D(_02975_),
    .Q(\cpuregs[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _26810_ (.CLK(clk),
    .D(_02976_),
    .Q(\cpuregs[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _26811_ (.CLK(clk),
    .D(_02977_),
    .Q(\cpuregs[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _26812_ (.CLK(clk),
    .D(_02978_),
    .Q(\cpuregs[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _26813_ (.CLK(clk),
    .D(_02979_),
    .Q(\cpuregs[2][16] ));
 sky130_fd_sc_hd__dfxtp_2 _26814_ (.CLK(clk),
    .D(_02980_),
    .Q(\cpuregs[2][17] ));
 sky130_fd_sc_hd__dfxtp_2 _26815_ (.CLK(clk),
    .D(_02981_),
    .Q(\cpuregs[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _26816_ (.CLK(clk),
    .D(_02982_),
    .Q(\cpuregs[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _26817_ (.CLK(clk),
    .D(_02983_),
    .Q(\cpuregs[2][20] ));
 sky130_fd_sc_hd__dfxtp_2 _26818_ (.CLK(clk),
    .D(_02984_),
    .Q(\cpuregs[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _26819_ (.CLK(clk),
    .D(_02985_),
    .Q(\cpuregs[2][22] ));
 sky130_fd_sc_hd__dfxtp_2 _26820_ (.CLK(clk),
    .D(_02986_),
    .Q(\cpuregs[2][23] ));
 sky130_fd_sc_hd__dfxtp_2 _26821_ (.CLK(clk),
    .D(_02987_),
    .Q(\cpuregs[2][24] ));
 sky130_fd_sc_hd__dfxtp_2 _26822_ (.CLK(clk),
    .D(_02988_),
    .Q(\cpuregs[2][25] ));
 sky130_fd_sc_hd__dfxtp_2 _26823_ (.CLK(clk),
    .D(_02989_),
    .Q(\cpuregs[2][26] ));
 sky130_fd_sc_hd__dfxtp_2 _26824_ (.CLK(clk),
    .D(_02990_),
    .Q(\cpuregs[2][27] ));
 sky130_fd_sc_hd__dfxtp_2 _26825_ (.CLK(clk),
    .D(_02991_),
    .Q(\cpuregs[2][28] ));
 sky130_fd_sc_hd__dfxtp_2 _26826_ (.CLK(clk),
    .D(_02992_),
    .Q(\cpuregs[2][29] ));
 sky130_fd_sc_hd__dfxtp_2 _26827_ (.CLK(clk),
    .D(_02993_),
    .Q(\cpuregs[2][30] ));
 sky130_fd_sc_hd__dfxtp_2 _26828_ (.CLK(clk),
    .D(_02994_),
    .Q(\cpuregs[2][31] ));
 sky130_fd_sc_hd__dfxtp_2 _26829_ (.CLK(clk),
    .D(_02995_),
    .Q(\cpuregs[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _26830_ (.CLK(clk),
    .D(_02996_),
    .Q(\cpuregs[5][1] ));
 sky130_fd_sc_hd__dfxtp_2 _26831_ (.CLK(clk),
    .D(_02997_),
    .Q(\cpuregs[5][2] ));
 sky130_fd_sc_hd__dfxtp_2 _26832_ (.CLK(clk),
    .D(_02998_),
    .Q(\cpuregs[5][3] ));
 sky130_fd_sc_hd__dfxtp_2 _26833_ (.CLK(clk),
    .D(_02999_),
    .Q(\cpuregs[5][4] ));
 sky130_fd_sc_hd__dfxtp_2 _26834_ (.CLK(clk),
    .D(_03000_),
    .Q(\cpuregs[5][5] ));
 sky130_fd_sc_hd__dfxtp_2 _26835_ (.CLK(clk),
    .D(_03001_),
    .Q(\cpuregs[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _26836_ (.CLK(clk),
    .D(_03002_),
    .Q(\cpuregs[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _26837_ (.CLK(clk),
    .D(_03003_),
    .Q(\cpuregs[5][8] ));
 sky130_fd_sc_hd__dfxtp_2 _26838_ (.CLK(clk),
    .D(_03004_),
    .Q(\cpuregs[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _26839_ (.CLK(clk),
    .D(_03005_),
    .Q(\cpuregs[5][10] ));
 sky130_fd_sc_hd__dfxtp_2 _26840_ (.CLK(clk),
    .D(_03006_),
    .Q(\cpuregs[5][11] ));
 sky130_fd_sc_hd__dfxtp_2 _26841_ (.CLK(clk),
    .D(_03007_),
    .Q(\cpuregs[5][12] ));
 sky130_fd_sc_hd__dfxtp_2 _26842_ (.CLK(clk),
    .D(_03008_),
    .Q(\cpuregs[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _26843_ (.CLK(clk),
    .D(_03009_),
    .Q(\cpuregs[5][14] ));
 sky130_fd_sc_hd__dfxtp_2 _26844_ (.CLK(clk),
    .D(_03010_),
    .Q(\cpuregs[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _26845_ (.CLK(clk),
    .D(_03011_),
    .Q(\cpuregs[5][16] ));
 sky130_fd_sc_hd__dfxtp_2 _26846_ (.CLK(clk),
    .D(_03012_),
    .Q(\cpuregs[5][17] ));
 sky130_fd_sc_hd__dfxtp_2 _26847_ (.CLK(clk),
    .D(_03013_),
    .Q(\cpuregs[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _26848_ (.CLK(clk),
    .D(_03014_),
    .Q(\cpuregs[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _26849_ (.CLK(clk),
    .D(_03015_),
    .Q(\cpuregs[5][20] ));
 sky130_fd_sc_hd__dfxtp_2 _26850_ (.CLK(clk),
    .D(_03016_),
    .Q(\cpuregs[5][21] ));
 sky130_fd_sc_hd__dfxtp_2 _26851_ (.CLK(clk),
    .D(_03017_),
    .Q(\cpuregs[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _26852_ (.CLK(clk),
    .D(_03018_),
    .Q(\cpuregs[5][23] ));
 sky130_fd_sc_hd__dfxtp_2 _26853_ (.CLK(clk),
    .D(_03019_),
    .Q(\cpuregs[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _26854_ (.CLK(clk),
    .D(_03020_),
    .Q(\cpuregs[5][25] ));
 sky130_fd_sc_hd__dfxtp_2 _26855_ (.CLK(clk),
    .D(_03021_),
    .Q(\cpuregs[5][26] ));
 sky130_fd_sc_hd__dfxtp_2 _26856_ (.CLK(clk),
    .D(_03022_),
    .Q(\cpuregs[5][27] ));
 sky130_fd_sc_hd__dfxtp_2 _26857_ (.CLK(clk),
    .D(_03023_),
    .Q(\cpuregs[5][28] ));
 sky130_fd_sc_hd__dfxtp_2 _26858_ (.CLK(clk),
    .D(_03024_),
    .Q(\cpuregs[5][29] ));
 sky130_fd_sc_hd__dfxtp_2 _26859_ (.CLK(clk),
    .D(_03025_),
    .Q(\cpuregs[5][30] ));
 sky130_fd_sc_hd__dfxtp_2 _26860_ (.CLK(clk),
    .D(_03026_),
    .Q(\cpuregs[5][31] ));
 sky130_fd_sc_hd__dfxtp_2 _26861_ (.CLK(clk),
    .D(_03027_),
    .Q(\pcpi_mul.rs1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _26862_ (.CLK(clk),
    .D(_03028_),
    .Q(\pcpi_mul.rs1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _26863_ (.CLK(clk),
    .D(_03029_),
    .Q(\pcpi_mul.rs1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _26864_ (.CLK(clk),
    .D(_03030_),
    .Q(\pcpi_mul.rs1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _26865_ (.CLK(clk),
    .D(_03031_),
    .Q(\pcpi_mul.rs1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _26866_ (.CLK(clk),
    .D(_03032_),
    .Q(\pcpi_mul.rs1[5] ));
 sky130_fd_sc_hd__dfxtp_2 _26867_ (.CLK(clk),
    .D(_03033_),
    .Q(\pcpi_mul.rs1[6] ));
 sky130_fd_sc_hd__dfxtp_2 _26868_ (.CLK(clk),
    .D(_03034_),
    .Q(\pcpi_mul.rs1[7] ));
 sky130_fd_sc_hd__dfxtp_2 _26869_ (.CLK(clk),
    .D(_03035_),
    .Q(\pcpi_mul.rs1[8] ));
 sky130_fd_sc_hd__dfxtp_2 _26870_ (.CLK(clk),
    .D(_03036_),
    .Q(\pcpi_mul.rs1[9] ));
 sky130_fd_sc_hd__dfxtp_2 _26871_ (.CLK(clk),
    .D(_03037_),
    .Q(\pcpi_mul.rs1[10] ));
 sky130_fd_sc_hd__dfxtp_2 _26872_ (.CLK(clk),
    .D(_03038_),
    .Q(\pcpi_mul.rs1[11] ));
 sky130_fd_sc_hd__dfxtp_2 _26873_ (.CLK(clk),
    .D(_03039_),
    .Q(\pcpi_mul.rs1[12] ));
 sky130_fd_sc_hd__dfxtp_2 _26874_ (.CLK(clk),
    .D(_03040_),
    .Q(\pcpi_mul.rs1[13] ));
 sky130_fd_sc_hd__dfxtp_2 _26875_ (.CLK(clk),
    .D(_03041_),
    .Q(\pcpi_mul.rs1[14] ));
 sky130_fd_sc_hd__dfxtp_2 _26876_ (.CLK(clk),
    .D(_03042_),
    .Q(\pcpi_mul.rs1[15] ));
 sky130_fd_sc_hd__dfxtp_2 _26877_ (.CLK(clk),
    .D(_03043_),
    .Q(\pcpi_mul.rs1[16] ));
 sky130_fd_sc_hd__dfxtp_2 _26878_ (.CLK(clk),
    .D(_03044_),
    .Q(\pcpi_mul.rs1[17] ));
 sky130_fd_sc_hd__dfxtp_2 _26879_ (.CLK(clk),
    .D(_03045_),
    .Q(\pcpi_mul.rs1[18] ));
 sky130_fd_sc_hd__dfxtp_2 _26880_ (.CLK(clk),
    .D(_03046_),
    .Q(\pcpi_mul.rs1[19] ));
 sky130_fd_sc_hd__dfxtp_2 _26881_ (.CLK(clk),
    .D(_03047_),
    .Q(\pcpi_mul.rs1[20] ));
 sky130_fd_sc_hd__dfxtp_2 _26882_ (.CLK(clk),
    .D(_03048_),
    .Q(\pcpi_mul.rs1[21] ));
 sky130_fd_sc_hd__dfxtp_2 _26883_ (.CLK(clk),
    .D(_03049_),
    .Q(\pcpi_mul.rs1[22] ));
 sky130_fd_sc_hd__dfxtp_2 _26884_ (.CLK(clk),
    .D(_03050_),
    .Q(\pcpi_mul.rs1[23] ));
 sky130_fd_sc_hd__dfxtp_2 _26885_ (.CLK(clk),
    .D(_03051_),
    .Q(\pcpi_mul.rs1[24] ));
 sky130_fd_sc_hd__dfxtp_2 _26886_ (.CLK(clk),
    .D(_03052_),
    .Q(\pcpi_mul.rs1[25] ));
 sky130_fd_sc_hd__dfxtp_2 _26887_ (.CLK(clk),
    .D(_03053_),
    .Q(\pcpi_mul.rs1[26] ));
 sky130_fd_sc_hd__dfxtp_2 _26888_ (.CLK(clk),
    .D(_03054_),
    .Q(\pcpi_mul.rs1[27] ));
 sky130_fd_sc_hd__dfxtp_2 _26889_ (.CLK(clk),
    .D(_03055_),
    .Q(\pcpi_mul.rs1[28] ));
 sky130_fd_sc_hd__dfxtp_2 _26890_ (.CLK(clk),
    .D(_03056_),
    .Q(\pcpi_mul.rs1[29] ));
 sky130_fd_sc_hd__dfxtp_2 _26891_ (.CLK(clk),
    .D(_03057_),
    .Q(\pcpi_mul.rs1[30] ));
 sky130_fd_sc_hd__dfxtp_2 _26892_ (.CLK(clk),
    .D(_03058_),
    .Q(\pcpi_mul.rs1[31] ));
 sky130_fd_sc_hd__dfxtp_2 _26893_ (.CLK(clk),
    .D(_03059_),
    .Q(mem_addr[2]));
 sky130_fd_sc_hd__dfxtp_2 _26894_ (.CLK(clk),
    .D(_03060_),
    .Q(mem_addr[3]));
 sky130_fd_sc_hd__dfxtp_2 _26895_ (.CLK(clk),
    .D(_03061_),
    .Q(mem_addr[4]));
 sky130_fd_sc_hd__dfxtp_2 _26896_ (.CLK(clk),
    .D(_03062_),
    .Q(mem_addr[5]));
 sky130_fd_sc_hd__dfxtp_2 _26897_ (.CLK(clk),
    .D(_03063_),
    .Q(mem_addr[6]));
 sky130_fd_sc_hd__dfxtp_2 _26898_ (.CLK(clk),
    .D(_03064_),
    .Q(mem_addr[7]));
 sky130_fd_sc_hd__dfxtp_2 _26899_ (.CLK(clk),
    .D(_03065_),
    .Q(mem_addr[8]));
 sky130_fd_sc_hd__dfxtp_2 _26900_ (.CLK(clk),
    .D(_03066_),
    .Q(mem_addr[9]));
 sky130_fd_sc_hd__dfxtp_2 _26901_ (.CLK(clk),
    .D(_03067_),
    .Q(mem_addr[10]));
 sky130_fd_sc_hd__dfxtp_2 _26902_ (.CLK(clk),
    .D(_03068_),
    .Q(mem_addr[11]));
 sky130_fd_sc_hd__dfxtp_2 _26903_ (.CLK(clk),
    .D(_03069_),
    .Q(mem_addr[12]));
 sky130_fd_sc_hd__dfxtp_2 _26904_ (.CLK(clk),
    .D(_03070_),
    .Q(mem_addr[13]));
 sky130_fd_sc_hd__dfxtp_2 _26905_ (.CLK(clk),
    .D(_03071_),
    .Q(mem_addr[14]));
 sky130_fd_sc_hd__dfxtp_2 _26906_ (.CLK(clk),
    .D(_03072_),
    .Q(mem_addr[15]));
 sky130_fd_sc_hd__dfxtp_2 _26907_ (.CLK(clk),
    .D(_03073_),
    .Q(mem_addr[16]));
 sky130_fd_sc_hd__dfxtp_2 _26908_ (.CLK(clk),
    .D(_03074_),
    .Q(mem_addr[17]));
 sky130_fd_sc_hd__dfxtp_2 _26909_ (.CLK(clk),
    .D(_03075_),
    .Q(mem_addr[18]));
 sky130_fd_sc_hd__dfxtp_2 _26910_ (.CLK(clk),
    .D(_03076_),
    .Q(mem_addr[19]));
 sky130_fd_sc_hd__dfxtp_2 _26911_ (.CLK(clk),
    .D(_03077_),
    .Q(mem_addr[20]));
 sky130_fd_sc_hd__dfxtp_2 _26912_ (.CLK(clk),
    .D(_03078_),
    .Q(mem_addr[21]));
 sky130_fd_sc_hd__dfxtp_2 _26913_ (.CLK(clk),
    .D(_03079_),
    .Q(mem_addr[22]));
 sky130_fd_sc_hd__dfxtp_2 _26914_ (.CLK(clk),
    .D(_03080_),
    .Q(mem_addr[23]));
 sky130_fd_sc_hd__dfxtp_2 _26915_ (.CLK(clk),
    .D(_03081_),
    .Q(mem_addr[24]));
 sky130_fd_sc_hd__dfxtp_2 _26916_ (.CLK(clk),
    .D(_03082_),
    .Q(mem_addr[25]));
 sky130_fd_sc_hd__dfxtp_2 _26917_ (.CLK(clk),
    .D(_03083_),
    .Q(mem_addr[26]));
 sky130_fd_sc_hd__dfxtp_2 _26918_ (.CLK(clk),
    .D(_03084_),
    .Q(mem_addr[27]));
 sky130_fd_sc_hd__dfxtp_2 _26919_ (.CLK(clk),
    .D(_03085_),
    .Q(mem_addr[28]));
 sky130_fd_sc_hd__dfxtp_2 _26920_ (.CLK(clk),
    .D(_03086_),
    .Q(mem_addr[29]));
 sky130_fd_sc_hd__dfxtp_2 _26921_ (.CLK(clk),
    .D(_03087_),
    .Q(mem_addr[30]));
 sky130_fd_sc_hd__dfxtp_2 _26922_ (.CLK(clk),
    .D(_03088_),
    .Q(mem_addr[31]));
 sky130_fd_sc_hd__dfxtp_2 _26923_ (.CLK(clk),
    .D(_03089_),
    .Q(pcpi_rs1[0]));
 sky130_fd_sc_hd__dfxtp_2 _26924_ (.CLK(clk),
    .D(_03090_),
    .Q(pcpi_rs1[1]));
 sky130_fd_sc_hd__dfxtp_2 _26925_ (.CLK(clk),
    .D(_03091_),
    .Q(pcpi_rs1[2]));
 sky130_fd_sc_hd__dfxtp_2 _26926_ (.CLK(clk),
    .D(_03092_),
    .Q(pcpi_rs1[3]));
 sky130_fd_sc_hd__dfxtp_2 _26927_ (.CLK(clk),
    .D(_03093_),
    .Q(pcpi_rs1[4]));
 sky130_fd_sc_hd__dfxtp_2 _26928_ (.CLK(clk),
    .D(_03094_),
    .Q(pcpi_rs1[5]));
 sky130_fd_sc_hd__dfxtp_2 _26929_ (.CLK(clk),
    .D(_03095_),
    .Q(pcpi_rs1[6]));
 sky130_fd_sc_hd__dfxtp_2 _26930_ (.CLK(clk),
    .D(_03096_),
    .Q(pcpi_rs1[7]));
 sky130_fd_sc_hd__dfxtp_2 _26931_ (.CLK(clk),
    .D(_03097_),
    .Q(pcpi_rs1[8]));
 sky130_fd_sc_hd__dfxtp_2 _26932_ (.CLK(clk),
    .D(_03098_),
    .Q(pcpi_rs1[9]));
 sky130_fd_sc_hd__dfxtp_2 _26933_ (.CLK(clk),
    .D(_03099_),
    .Q(pcpi_rs1[10]));
 sky130_fd_sc_hd__dfxtp_2 _26934_ (.CLK(clk),
    .D(_03100_),
    .Q(pcpi_rs1[11]));
 sky130_fd_sc_hd__dfxtp_2 _26935_ (.CLK(clk),
    .D(_03101_),
    .Q(pcpi_rs1[12]));
 sky130_fd_sc_hd__dfxtp_2 _26936_ (.CLK(clk),
    .D(_03102_),
    .Q(pcpi_rs1[13]));
 sky130_fd_sc_hd__dfxtp_2 _26937_ (.CLK(clk),
    .D(_03103_),
    .Q(pcpi_rs1[14]));
 sky130_fd_sc_hd__dfxtp_2 _26938_ (.CLK(clk),
    .D(_03104_),
    .Q(pcpi_rs1[15]));
 sky130_fd_sc_hd__dfxtp_2 _26939_ (.CLK(clk),
    .D(_03105_),
    .Q(pcpi_rs1[16]));
 sky130_fd_sc_hd__dfxtp_2 _26940_ (.CLK(clk),
    .D(_03106_),
    .Q(pcpi_rs1[17]));
 sky130_fd_sc_hd__dfxtp_2 _26941_ (.CLK(clk),
    .D(_03107_),
    .Q(pcpi_rs1[18]));
 sky130_fd_sc_hd__dfxtp_2 _26942_ (.CLK(clk),
    .D(_03108_),
    .Q(pcpi_rs1[19]));
 sky130_fd_sc_hd__dfxtp_2 _26943_ (.CLK(clk),
    .D(_03109_),
    .Q(pcpi_rs1[20]));
 sky130_fd_sc_hd__dfxtp_2 _26944_ (.CLK(clk),
    .D(_03110_),
    .Q(pcpi_rs1[21]));
 sky130_fd_sc_hd__dfxtp_2 _26945_ (.CLK(clk),
    .D(_03111_),
    .Q(pcpi_rs1[22]));
 sky130_fd_sc_hd__dfxtp_2 _26946_ (.CLK(clk),
    .D(_03112_),
    .Q(pcpi_rs1[23]));
 sky130_fd_sc_hd__dfxtp_2 _26947_ (.CLK(clk),
    .D(_03113_),
    .Q(pcpi_rs1[24]));
 sky130_fd_sc_hd__dfxtp_2 _26948_ (.CLK(clk),
    .D(_03114_),
    .Q(pcpi_rs1[25]));
 sky130_fd_sc_hd__dfxtp_2 _26949_ (.CLK(clk),
    .D(_03115_),
    .Q(pcpi_rs1[26]));
 sky130_fd_sc_hd__dfxtp_2 _26950_ (.CLK(clk),
    .D(_03116_),
    .Q(pcpi_rs1[27]));
 sky130_fd_sc_hd__dfxtp_2 _26951_ (.CLK(clk),
    .D(_03117_),
    .Q(pcpi_rs1[28]));
 sky130_fd_sc_hd__dfxtp_2 _26952_ (.CLK(clk),
    .D(_03118_),
    .Q(pcpi_rs1[29]));
 sky130_fd_sc_hd__dfxtp_2 _26953_ (.CLK(clk),
    .D(_03119_),
    .Q(pcpi_rs1[30]));
 sky130_fd_sc_hd__dfxtp_2 _26954_ (.CLK(clk),
    .D(_03120_),
    .Q(pcpi_rs1[31]));
 sky130_fd_sc_hd__dfxtp_2 _26955_ (.CLK(clk),
    .D(_03121_),
    .Q(pcpi_insn[0]));
 sky130_fd_sc_hd__dfxtp_2 _26956_ (.CLK(clk),
    .D(_03122_),
    .Q(pcpi_insn[1]));
 sky130_fd_sc_hd__dfxtp_2 _26957_ (.CLK(clk),
    .D(_03123_),
    .Q(pcpi_insn[2]));
 sky130_fd_sc_hd__dfxtp_2 _26958_ (.CLK(clk),
    .D(_03124_),
    .Q(pcpi_insn[3]));
 sky130_fd_sc_hd__dfxtp_2 _26959_ (.CLK(clk),
    .D(_03125_),
    .Q(pcpi_insn[4]));
 sky130_fd_sc_hd__dfxtp_2 _26960_ (.CLK(clk),
    .D(_03126_),
    .Q(pcpi_insn[5]));
 sky130_fd_sc_hd__dfxtp_2 _26961_ (.CLK(clk),
    .D(_03127_),
    .Q(pcpi_insn[6]));
 sky130_fd_sc_hd__dfxtp_2 _26962_ (.CLK(clk),
    .D(_03128_),
    .Q(pcpi_insn[7]));
 sky130_fd_sc_hd__dfxtp_2 _26963_ (.CLK(clk),
    .D(_03129_),
    .Q(pcpi_insn[8]));
 sky130_fd_sc_hd__dfxtp_2 _26964_ (.CLK(clk),
    .D(_03130_),
    .Q(pcpi_insn[9]));
 sky130_fd_sc_hd__dfxtp_2 _26965_ (.CLK(clk),
    .D(_03131_),
    .Q(pcpi_insn[10]));
 sky130_fd_sc_hd__dfxtp_2 _26966_ (.CLK(clk),
    .D(_03132_),
    .Q(pcpi_insn[11]));
 sky130_fd_sc_hd__dfxtp_2 _26967_ (.CLK(clk),
    .D(_03133_),
    .Q(pcpi_insn[12]));
 sky130_fd_sc_hd__dfxtp_2 _26968_ (.CLK(clk),
    .D(_03134_),
    .Q(pcpi_insn[13]));
 sky130_fd_sc_hd__dfxtp_2 _26969_ (.CLK(clk),
    .D(_03135_),
    .Q(pcpi_insn[14]));
 sky130_fd_sc_hd__dfxtp_2 _26970_ (.CLK(clk),
    .D(_03136_),
    .Q(pcpi_insn[15]));
 sky130_fd_sc_hd__dfxtp_2 _26971_ (.CLK(clk),
    .D(_03137_),
    .Q(pcpi_insn[16]));
 sky130_fd_sc_hd__dfxtp_2 _26972_ (.CLK(clk),
    .D(_03138_),
    .Q(pcpi_insn[17]));
 sky130_fd_sc_hd__dfxtp_2 _26973_ (.CLK(clk),
    .D(_03139_),
    .Q(pcpi_insn[18]));
 sky130_fd_sc_hd__dfxtp_2 _26974_ (.CLK(clk),
    .D(_03140_),
    .Q(pcpi_insn[19]));
 sky130_fd_sc_hd__dfxtp_2 _26975_ (.CLK(clk),
    .D(_03141_),
    .Q(pcpi_insn[20]));
 sky130_fd_sc_hd__dfxtp_2 _26976_ (.CLK(clk),
    .D(_03142_),
    .Q(pcpi_insn[21]));
 sky130_fd_sc_hd__dfxtp_2 _26977_ (.CLK(clk),
    .D(_03143_),
    .Q(pcpi_insn[22]));
 sky130_fd_sc_hd__dfxtp_2 _26978_ (.CLK(clk),
    .D(_03144_),
    .Q(pcpi_insn[23]));
 sky130_fd_sc_hd__dfxtp_2 _26979_ (.CLK(clk),
    .D(_03145_),
    .Q(pcpi_insn[24]));
 sky130_fd_sc_hd__dfxtp_2 _26980_ (.CLK(clk),
    .D(_03146_),
    .Q(pcpi_insn[25]));
 sky130_fd_sc_hd__dfxtp_2 _26981_ (.CLK(clk),
    .D(_03147_),
    .Q(pcpi_insn[26]));
 sky130_fd_sc_hd__dfxtp_2 _26982_ (.CLK(clk),
    .D(_03148_),
    .Q(pcpi_insn[27]));
 sky130_fd_sc_hd__dfxtp_2 _26983_ (.CLK(clk),
    .D(_03149_),
    .Q(pcpi_insn[28]));
 sky130_fd_sc_hd__dfxtp_2 _26984_ (.CLK(clk),
    .D(_03150_),
    .Q(pcpi_insn[29]));
 sky130_fd_sc_hd__dfxtp_2 _26985_ (.CLK(clk),
    .D(_03151_),
    .Q(pcpi_insn[30]));
 sky130_fd_sc_hd__dfxtp_2 _26986_ (.CLK(clk),
    .D(_03152_),
    .Q(pcpi_insn[31]));
 sky130_fd_sc_hd__dfxtp_2 _26987_ (.CLK(clk),
    .D(_03153_),
    .Q(instr_lui));
 sky130_fd_sc_hd__dfxtp_2 _26988_ (.CLK(clk),
    .D(_03154_),
    .Q(instr_auipc));
 sky130_fd_sc_hd__dfxtp_2 _26989_ (.CLK(clk),
    .D(_03155_),
    .Q(instr_jal));
 sky130_fd_sc_hd__dfxtp_2 _26990_ (.CLK(clk),
    .D(_03156_),
    .Q(instr_jalr));
 sky130_fd_sc_hd__dfxtp_2 _26991_ (.CLK(clk),
    .D(_03157_),
    .Q(instr_lb));
 sky130_fd_sc_hd__dfxtp_2 _26992_ (.CLK(clk),
    .D(_03158_),
    .Q(instr_lh));
 sky130_fd_sc_hd__dfxtp_2 _26993_ (.CLK(clk),
    .D(_03159_),
    .Q(instr_lw));
 sky130_fd_sc_hd__dfxtp_2 _26994_ (.CLK(clk),
    .D(_03160_),
    .Q(instr_lbu));
 sky130_fd_sc_hd__dfxtp_2 _26995_ (.CLK(clk),
    .D(_03161_),
    .Q(instr_lhu));
 sky130_fd_sc_hd__dfxtp_2 _26996_ (.CLK(clk),
    .D(_03162_),
    .Q(instr_sb));
 sky130_fd_sc_hd__dfxtp_2 _26997_ (.CLK(clk),
    .D(_03163_),
    .Q(instr_sh));
 sky130_fd_sc_hd__dfxtp_2 _26998_ (.CLK(clk),
    .D(_03164_),
    .Q(instr_sw));
 sky130_fd_sc_hd__dfxtp_2 _26999_ (.CLK(clk),
    .D(_03165_),
    .Q(instr_slli));
 sky130_fd_sc_hd__dfxtp_2 _27000_ (.CLK(clk),
    .D(_03166_),
    .Q(instr_srli));
 sky130_fd_sc_hd__dfxtp_2 _27001_ (.CLK(clk),
    .D(_03167_),
    .Q(instr_srai));
 sky130_fd_sc_hd__dfxtp_2 _27002_ (.CLK(clk),
    .D(_03168_),
    .Q(instr_rdcycle));
 sky130_fd_sc_hd__dfxtp_2 _27003_ (.CLK(clk),
    .D(_03169_),
    .Q(instr_rdcycleh));
 sky130_fd_sc_hd__dfxtp_2 _27004_ (.CLK(clk),
    .D(_03170_),
    .Q(instr_rdinstr));
 sky130_fd_sc_hd__dfxtp_2 _27005_ (.CLK(clk),
    .D(_03171_),
    .Q(instr_rdinstrh));
 sky130_fd_sc_hd__dfxtp_2 _27006_ (.CLK(clk),
    .D(_03172_),
    .Q(instr_ecall_ebreak));
 sky130_fd_sc_hd__dfxtp_2 _27007_ (.CLK(clk),
    .D(_03173_),
    .Q(instr_getq));
 sky130_fd_sc_hd__dfxtp_2 _27008_ (.CLK(clk),
    .D(_03174_),
    .Q(instr_setq));
 sky130_fd_sc_hd__dfxtp_2 _27009_ (.CLK(clk),
    .D(_03175_),
    .Q(instr_retirq));
 sky130_fd_sc_hd__dfxtp_2 _27010_ (.CLK(clk),
    .D(_03176_),
    .Q(instr_maskirq));
 sky130_fd_sc_hd__dfxtp_2 _27011_ (.CLK(clk),
    .D(_03177_),
    .Q(instr_waitirq));
 sky130_fd_sc_hd__dfxtp_2 _27012_ (.CLK(clk),
    .D(_03178_),
    .Q(instr_timer));
 sky130_fd_sc_hd__dfxtp_2 _27013_ (.CLK(clk),
    .D(_03179_),
    .Q(\decoded_rd[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27014_ (.CLK(clk),
    .D(_03180_),
    .Q(\decoded_rd[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27015_ (.CLK(clk),
    .D(_03181_),
    .Q(\decoded_rd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27016_ (.CLK(clk),
    .D(_03182_),
    .Q(\decoded_rd[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27017_ (.CLK(clk),
    .D(_03183_),
    .Q(\decoded_rd[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27018_ (.CLK(clk),
    .D(_03184_),
    .Q(\decoded_imm[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27019_ (.CLK(clk),
    .D(_03185_),
    .Q(\decoded_imm_uj[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27020_ (.CLK(clk),
    .D(_03186_),
    .Q(\decoded_imm_uj[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27021_ (.CLK(clk),
    .D(_03187_),
    .Q(\decoded_imm_uj[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27022_ (.CLK(clk),
    .D(_03188_),
    .Q(\decoded_imm_uj[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27023_ (.CLK(clk),
    .D(_03189_),
    .Q(\decoded_imm_uj[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27024_ (.CLK(clk),
    .D(_03190_),
    .Q(\decoded_imm_uj[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27025_ (.CLK(clk),
    .D(_03191_),
    .Q(\decoded_imm_uj[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27026_ (.CLK(clk),
    .D(_03192_),
    .Q(\decoded_imm_uj[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27027_ (.CLK(clk),
    .D(_03193_),
    .Q(\decoded_imm_uj[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27028_ (.CLK(clk),
    .D(_03194_),
    .Q(\decoded_imm_uj[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27029_ (.CLK(clk),
    .D(_03195_),
    .Q(\decoded_imm_uj[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27030_ (.CLK(clk),
    .D(_03196_),
    .Q(\decoded_imm_uj[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27031_ (.CLK(clk),
    .D(_03197_),
    .Q(\decoded_imm_uj[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27032_ (.CLK(clk),
    .D(_03198_),
    .Q(\decoded_imm_uj[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27033_ (.CLK(clk),
    .D(_03199_),
    .Q(\decoded_imm_uj[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27034_ (.CLK(clk),
    .D(_03200_),
    .Q(\decoded_imm_uj[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27035_ (.CLK(clk),
    .D(_03201_),
    .Q(\decoded_imm_uj[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27036_ (.CLK(clk),
    .D(_03202_),
    .Q(\decoded_imm_uj[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27037_ (.CLK(clk),
    .D(_03203_),
    .Q(\decoded_imm_uj[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27038_ (.CLK(clk),
    .D(_03204_),
    .Q(\decoded_imm_uj[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27039_ (.CLK(clk),
    .D(_03205_),
    .Q(is_lb_lh_lw_lbu_lhu));
 sky130_fd_sc_hd__dfxtp_2 _27040_ (.CLK(clk),
    .D(_03206_),
    .Q(is_slli_srli_srai));
 sky130_fd_sc_hd__dfxtp_2 _27041_ (.CLK(clk),
    .D(_03207_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi));
 sky130_fd_sc_hd__dfxtp_2 _27042_ (.CLK(clk),
    .D(_03208_),
    .Q(is_sb_sh_sw));
 sky130_fd_sc_hd__dfxtp_2 _27043_ (.CLK(clk),
    .D(_03209_),
    .Q(\cpuregs[13][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27044_ (.CLK(clk),
    .D(_03210_),
    .Q(\cpuregs[13][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27045_ (.CLK(clk),
    .D(_03211_),
    .Q(\cpuregs[13][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27046_ (.CLK(clk),
    .D(_03212_),
    .Q(\cpuregs[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27047_ (.CLK(clk),
    .D(_03213_),
    .Q(\cpuregs[13][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27048_ (.CLK(clk),
    .D(_03214_),
    .Q(\cpuregs[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27049_ (.CLK(clk),
    .D(_03215_),
    .Q(\cpuregs[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27050_ (.CLK(clk),
    .D(_03216_),
    .Q(\cpuregs[13][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27051_ (.CLK(clk),
    .D(_03217_),
    .Q(\cpuregs[13][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27052_ (.CLK(clk),
    .D(_03218_),
    .Q(\cpuregs[13][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27053_ (.CLK(clk),
    .D(_03219_),
    .Q(\cpuregs[13][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27054_ (.CLK(clk),
    .D(_03220_),
    .Q(\cpuregs[13][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27055_ (.CLK(clk),
    .D(_03221_),
    .Q(\cpuregs[13][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27056_ (.CLK(clk),
    .D(_03222_),
    .Q(\cpuregs[13][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27057_ (.CLK(clk),
    .D(_03223_),
    .Q(\cpuregs[13][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27058_ (.CLK(clk),
    .D(_03224_),
    .Q(\cpuregs[13][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27059_ (.CLK(clk),
    .D(_03225_),
    .Q(\cpuregs[13][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27060_ (.CLK(clk),
    .D(_03226_),
    .Q(\cpuregs[13][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27061_ (.CLK(clk),
    .D(_03227_),
    .Q(\cpuregs[13][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27062_ (.CLK(clk),
    .D(_03228_),
    .Q(\cpuregs[13][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27063_ (.CLK(clk),
    .D(_03229_),
    .Q(\cpuregs[13][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27064_ (.CLK(clk),
    .D(_03230_),
    .Q(\cpuregs[13][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27065_ (.CLK(clk),
    .D(_03231_),
    .Q(\cpuregs[13][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27066_ (.CLK(clk),
    .D(_03232_),
    .Q(\cpuregs[13][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27067_ (.CLK(clk),
    .D(_03233_),
    .Q(\cpuregs[13][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27068_ (.CLK(clk),
    .D(_03234_),
    .Q(\cpuregs[13][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27069_ (.CLK(clk),
    .D(_03235_),
    .Q(\cpuregs[13][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27070_ (.CLK(clk),
    .D(_03236_),
    .Q(\cpuregs[13][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27071_ (.CLK(clk),
    .D(_03237_),
    .Q(\cpuregs[13][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27072_ (.CLK(clk),
    .D(_03238_),
    .Q(\cpuregs[13][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27073_ (.CLK(clk),
    .D(_03239_),
    .Q(\cpuregs[13][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27074_ (.CLK(clk),
    .D(_03240_),
    .Q(\cpuregs[13][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27075_ (.CLK(clk),
    .D(_03241_),
    .Q(is_alu_reg_imm));
 sky130_fd_sc_hd__dfxtp_2 _27076_ (.CLK(clk),
    .D(_03242_),
    .Q(is_alu_reg_reg));
 sky130_fd_sc_hd__dfxtp_2 _27077_ (.CLK(clk),
    .D(_03243_),
    .Q(mem_wstrb[0]));
 sky130_fd_sc_hd__dfxtp_2 _27078_ (.CLK(clk),
    .D(_03244_),
    .Q(mem_wstrb[1]));
 sky130_fd_sc_hd__dfxtp_2 _27079_ (.CLK(clk),
    .D(_03245_),
    .Q(mem_wstrb[2]));
 sky130_fd_sc_hd__dfxtp_2 _27080_ (.CLK(clk),
    .D(_03246_),
    .Q(mem_wstrb[3]));
 sky130_fd_sc_hd__dfxtp_2 _27081_ (.CLK(clk),
    .D(_03247_),
    .Q(\pcpi_mul.rs2[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27082_ (.CLK(clk),
    .D(_03248_),
    .Q(\pcpi_mul.rs2[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27083_ (.CLK(clk),
    .D(_03249_),
    .Q(\pcpi_mul.rs2[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27084_ (.CLK(clk),
    .D(_03250_),
    .Q(\pcpi_mul.rs2[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27085_ (.CLK(clk),
    .D(_03251_),
    .Q(\pcpi_mul.rs2[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27086_ (.CLK(clk),
    .D(_03252_),
    .Q(\pcpi_mul.rs2[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27087_ (.CLK(clk),
    .D(_03253_),
    .Q(\pcpi_mul.rs2[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27088_ (.CLK(clk),
    .D(_03254_),
    .Q(\pcpi_mul.rs2[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27089_ (.CLK(clk),
    .D(_03255_),
    .Q(\pcpi_mul.rs2[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27090_ (.CLK(clk),
    .D(_03256_),
    .Q(\pcpi_mul.rs2[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27091_ (.CLK(clk),
    .D(_03257_),
    .Q(\pcpi_mul.rs2[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27092_ (.CLK(clk),
    .D(_03258_),
    .Q(\pcpi_mul.rs2[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27093_ (.CLK(clk),
    .D(_03259_),
    .Q(\pcpi_mul.rs2[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27094_ (.CLK(clk),
    .D(_03260_),
    .Q(\pcpi_mul.rs2[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27095_ (.CLK(clk),
    .D(_03261_),
    .Q(\pcpi_mul.rs2[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27096_ (.CLK(clk),
    .D(_03262_),
    .Q(\pcpi_mul.rs2[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27097_ (.CLK(clk),
    .D(_03263_),
    .Q(\pcpi_mul.rs2[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27098_ (.CLK(clk),
    .D(_03264_),
    .Q(\pcpi_mul.rs2[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27099_ (.CLK(clk),
    .D(_03265_),
    .Q(\pcpi_mul.rs2[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27100_ (.CLK(clk),
    .D(_03266_),
    .Q(\pcpi_mul.rs2[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27101_ (.CLK(clk),
    .D(_03267_),
    .Q(\pcpi_mul.rs2[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27102_ (.CLK(clk),
    .D(_03268_),
    .Q(\pcpi_mul.rs2[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27103_ (.CLK(clk),
    .D(_03269_),
    .Q(\pcpi_mul.rs2[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27104_ (.CLK(clk),
    .D(_03270_),
    .Q(\pcpi_mul.rs2[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27105_ (.CLK(clk),
    .D(_03271_),
    .Q(\pcpi_mul.rs2[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27106_ (.CLK(clk),
    .D(_03272_),
    .Q(\pcpi_mul.rs2[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27107_ (.CLK(clk),
    .D(_03273_),
    .Q(\pcpi_mul.rs2[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27108_ (.CLK(clk),
    .D(_03274_),
    .Q(\pcpi_mul.rs2[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27109_ (.CLK(clk),
    .D(_03275_),
    .Q(\pcpi_mul.rs2[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27110_ (.CLK(clk),
    .D(_03276_),
    .Q(\pcpi_mul.rs2[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27111_ (.CLK(clk),
    .D(_03277_),
    .Q(\pcpi_mul.rs2[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27112_ (.CLK(clk),
    .D(_03278_),
    .Q(\pcpi_mul.rs2[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27113_ (.CLK(clk),
    .D(_03279_),
    .Q(\cpuregs[17][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27114_ (.CLK(clk),
    .D(_03280_),
    .Q(\cpuregs[17][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27115_ (.CLK(clk),
    .D(_03281_),
    .Q(\cpuregs[17][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27116_ (.CLK(clk),
    .D(_03282_),
    .Q(\cpuregs[17][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27117_ (.CLK(clk),
    .D(_03283_),
    .Q(\cpuregs[17][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27118_ (.CLK(clk),
    .D(_03284_),
    .Q(\cpuregs[17][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27119_ (.CLK(clk),
    .D(_03285_),
    .Q(\cpuregs[17][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27120_ (.CLK(clk),
    .D(_03286_),
    .Q(\cpuregs[17][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27121_ (.CLK(clk),
    .D(_03287_),
    .Q(\cpuregs[17][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27122_ (.CLK(clk),
    .D(_03288_),
    .Q(\cpuregs[17][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27123_ (.CLK(clk),
    .D(_03289_),
    .Q(\cpuregs[17][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27124_ (.CLK(clk),
    .D(_03290_),
    .Q(\cpuregs[17][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27125_ (.CLK(clk),
    .D(_03291_),
    .Q(\cpuregs[17][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27126_ (.CLK(clk),
    .D(_03292_),
    .Q(\cpuregs[17][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27127_ (.CLK(clk),
    .D(_03293_),
    .Q(\cpuregs[17][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27128_ (.CLK(clk),
    .D(_03294_),
    .Q(\cpuregs[17][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27129_ (.CLK(clk),
    .D(_03295_),
    .Q(\cpuregs[17][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27130_ (.CLK(clk),
    .D(_03296_),
    .Q(\cpuregs[17][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27131_ (.CLK(clk),
    .D(_03297_),
    .Q(\cpuregs[17][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27132_ (.CLK(clk),
    .D(_03298_),
    .Q(\cpuregs[17][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27133_ (.CLK(clk),
    .D(_03299_),
    .Q(\cpuregs[17][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27134_ (.CLK(clk),
    .D(_03300_),
    .Q(\cpuregs[17][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27135_ (.CLK(clk),
    .D(_03301_),
    .Q(\cpuregs[17][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27136_ (.CLK(clk),
    .D(_03302_),
    .Q(\cpuregs[17][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27137_ (.CLK(clk),
    .D(_03303_),
    .Q(\cpuregs[17][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27138_ (.CLK(clk),
    .D(_03304_),
    .Q(\cpuregs[17][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27139_ (.CLK(clk),
    .D(_03305_),
    .Q(\cpuregs[17][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27140_ (.CLK(clk),
    .D(_03306_),
    .Q(\cpuregs[17][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27141_ (.CLK(clk),
    .D(_03307_),
    .Q(\cpuregs[17][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27142_ (.CLK(clk),
    .D(_03308_),
    .Q(\cpuregs[17][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27143_ (.CLK(clk),
    .D(_03309_),
    .Q(\cpuregs[17][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27144_ (.CLK(clk),
    .D(_03310_),
    .Q(\cpuregs[17][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27145_ (.CLK(clk),
    .D(_03311_),
    .Q(\cpuregs[16][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27146_ (.CLK(clk),
    .D(_03312_),
    .Q(\cpuregs[16][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27147_ (.CLK(clk),
    .D(_03313_),
    .Q(\cpuregs[16][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27148_ (.CLK(clk),
    .D(_03314_),
    .Q(\cpuregs[16][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27149_ (.CLK(clk),
    .D(_03315_),
    .Q(\cpuregs[16][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27150_ (.CLK(clk),
    .D(_03316_),
    .Q(\cpuregs[16][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27151_ (.CLK(clk),
    .D(_03317_),
    .Q(\cpuregs[16][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27152_ (.CLK(clk),
    .D(_03318_),
    .Q(\cpuregs[16][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27153_ (.CLK(clk),
    .D(_03319_),
    .Q(\cpuregs[16][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27154_ (.CLK(clk),
    .D(_03320_),
    .Q(\cpuregs[16][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27155_ (.CLK(clk),
    .D(_03321_),
    .Q(\cpuregs[16][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27156_ (.CLK(clk),
    .D(_03322_),
    .Q(\cpuregs[16][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27157_ (.CLK(clk),
    .D(_03323_),
    .Q(\cpuregs[16][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27158_ (.CLK(clk),
    .D(_03324_),
    .Q(\cpuregs[16][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27159_ (.CLK(clk),
    .D(_03325_),
    .Q(\cpuregs[16][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27160_ (.CLK(clk),
    .D(_03326_),
    .Q(\cpuregs[16][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27161_ (.CLK(clk),
    .D(_03327_),
    .Q(\cpuregs[16][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27162_ (.CLK(clk),
    .D(_03328_),
    .Q(\cpuregs[16][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27163_ (.CLK(clk),
    .D(_03329_),
    .Q(\cpuregs[16][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27164_ (.CLK(clk),
    .D(_03330_),
    .Q(\cpuregs[16][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27165_ (.CLK(clk),
    .D(_03331_),
    .Q(\cpuregs[16][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27166_ (.CLK(clk),
    .D(_03332_),
    .Q(\cpuregs[16][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27167_ (.CLK(clk),
    .D(_03333_),
    .Q(\cpuregs[16][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27168_ (.CLK(clk),
    .D(_03334_),
    .Q(\cpuregs[16][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27169_ (.CLK(clk),
    .D(_03335_),
    .Q(\cpuregs[16][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27170_ (.CLK(clk),
    .D(_03336_),
    .Q(\cpuregs[16][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27171_ (.CLK(clk),
    .D(_03337_),
    .Q(\cpuregs[16][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27172_ (.CLK(clk),
    .D(_03338_),
    .Q(\cpuregs[16][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27173_ (.CLK(clk),
    .D(_03339_),
    .Q(\cpuregs[16][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27174_ (.CLK(clk),
    .D(_03340_),
    .Q(\cpuregs[16][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27175_ (.CLK(clk),
    .D(_03341_),
    .Q(\cpuregs[16][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27176_ (.CLK(clk),
    .D(_03342_),
    .Q(\cpuregs[16][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27177_ (.CLK(clk),
    .D(_03343_),
    .Q(\cpuregs[12][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27178_ (.CLK(clk),
    .D(_03344_),
    .Q(\cpuregs[12][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27179_ (.CLK(clk),
    .D(_03345_),
    .Q(\cpuregs[12][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27180_ (.CLK(clk),
    .D(_03346_),
    .Q(\cpuregs[12][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27181_ (.CLK(clk),
    .D(_03347_),
    .Q(\cpuregs[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27182_ (.CLK(clk),
    .D(_03348_),
    .Q(\cpuregs[12][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27183_ (.CLK(clk),
    .D(_03349_),
    .Q(\cpuregs[12][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27184_ (.CLK(clk),
    .D(_03350_),
    .Q(\cpuregs[12][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27185_ (.CLK(clk),
    .D(_03351_),
    .Q(\cpuregs[12][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27186_ (.CLK(clk),
    .D(_03352_),
    .Q(\cpuregs[12][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27187_ (.CLK(clk),
    .D(_03353_),
    .Q(\cpuregs[12][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27188_ (.CLK(clk),
    .D(_03354_),
    .Q(\cpuregs[12][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27189_ (.CLK(clk),
    .D(_03355_),
    .Q(\cpuregs[12][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27190_ (.CLK(clk),
    .D(_03356_),
    .Q(\cpuregs[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27191_ (.CLK(clk),
    .D(_03357_),
    .Q(\cpuregs[12][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27192_ (.CLK(clk),
    .D(_03358_),
    .Q(\cpuregs[12][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27193_ (.CLK(clk),
    .D(_03359_),
    .Q(\cpuregs[12][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27194_ (.CLK(clk),
    .D(_03360_),
    .Q(\cpuregs[12][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27195_ (.CLK(clk),
    .D(_03361_),
    .Q(\cpuregs[12][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27196_ (.CLK(clk),
    .D(_03362_),
    .Q(\cpuregs[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27197_ (.CLK(clk),
    .D(_03363_),
    .Q(\cpuregs[12][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27198_ (.CLK(clk),
    .D(_03364_),
    .Q(\cpuregs[12][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27199_ (.CLK(clk),
    .D(_03365_),
    .Q(\cpuregs[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27200_ (.CLK(clk),
    .D(_03366_),
    .Q(\cpuregs[12][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27201_ (.CLK(clk),
    .D(_03367_),
    .Q(\cpuregs[12][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27202_ (.CLK(clk),
    .D(_03368_),
    .Q(\cpuregs[12][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27203_ (.CLK(clk),
    .D(_03369_),
    .Q(\cpuregs[12][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27204_ (.CLK(clk),
    .D(_03370_),
    .Q(\cpuregs[12][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27205_ (.CLK(clk),
    .D(_03371_),
    .Q(\cpuregs[12][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27206_ (.CLK(clk),
    .D(_03372_),
    .Q(\cpuregs[12][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27207_ (.CLK(clk),
    .D(_03373_),
    .Q(\cpuregs[12][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27208_ (.CLK(clk),
    .D(_03374_),
    .Q(\cpuregs[12][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27209_ (.CLK(clk),
    .D(_03375_),
    .Q(\cpuregs[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27210_ (.CLK(clk),
    .D(_03376_),
    .Q(\cpuregs[1][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27211_ (.CLK(clk),
    .D(_03377_),
    .Q(\cpuregs[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27212_ (.CLK(clk),
    .D(_03378_),
    .Q(\cpuregs[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27213_ (.CLK(clk),
    .D(_03379_),
    .Q(\cpuregs[1][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27214_ (.CLK(clk),
    .D(_03380_),
    .Q(\cpuregs[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27215_ (.CLK(clk),
    .D(_03381_),
    .Q(\cpuregs[1][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27216_ (.CLK(clk),
    .D(_03382_),
    .Q(\cpuregs[1][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27217_ (.CLK(clk),
    .D(_03383_),
    .Q(\cpuregs[1][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27218_ (.CLK(clk),
    .D(_03384_),
    .Q(\cpuregs[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27219_ (.CLK(clk),
    .D(_03385_),
    .Q(\cpuregs[1][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27220_ (.CLK(clk),
    .D(_03386_),
    .Q(\cpuregs[1][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27221_ (.CLK(clk),
    .D(_03387_),
    .Q(\cpuregs[1][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27222_ (.CLK(clk),
    .D(_03388_),
    .Q(\cpuregs[1][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27223_ (.CLK(clk),
    .D(_03389_),
    .Q(\cpuregs[1][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27224_ (.CLK(clk),
    .D(_03390_),
    .Q(\cpuregs[1][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27225_ (.CLK(clk),
    .D(_03391_),
    .Q(\cpuregs[1][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27226_ (.CLK(clk),
    .D(_03392_),
    .Q(\cpuregs[1][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27227_ (.CLK(clk),
    .D(_03393_),
    .Q(\cpuregs[1][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27228_ (.CLK(clk),
    .D(_03394_),
    .Q(\cpuregs[1][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27229_ (.CLK(clk),
    .D(_03395_),
    .Q(\cpuregs[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27230_ (.CLK(clk),
    .D(_03396_),
    .Q(\cpuregs[1][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27231_ (.CLK(clk),
    .D(_03397_),
    .Q(\cpuregs[1][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27232_ (.CLK(clk),
    .D(_03398_),
    .Q(\cpuregs[1][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27233_ (.CLK(clk),
    .D(_03399_),
    .Q(\cpuregs[1][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27234_ (.CLK(clk),
    .D(_03400_),
    .Q(\cpuregs[1][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27235_ (.CLK(clk),
    .D(_03401_),
    .Q(\cpuregs[1][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27236_ (.CLK(clk),
    .D(_03402_),
    .Q(\cpuregs[1][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27237_ (.CLK(clk),
    .D(_03403_),
    .Q(\cpuregs[1][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27238_ (.CLK(clk),
    .D(_03404_),
    .Q(\cpuregs[1][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27239_ (.CLK(clk),
    .D(_03405_),
    .Q(\cpuregs[1][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27240_ (.CLK(clk),
    .D(_03406_),
    .Q(\cpuregs[1][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27241_ (.CLK(clk),
    .D(_03407_),
    .Q(\cpuregs[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27242_ (.CLK(clk),
    .D(_03408_),
    .Q(\cpuregs[3][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27243_ (.CLK(clk),
    .D(_03409_),
    .Q(\cpuregs[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27244_ (.CLK(clk),
    .D(_03410_),
    .Q(\cpuregs[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27245_ (.CLK(clk),
    .D(_03411_),
    .Q(\cpuregs[3][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27246_ (.CLK(clk),
    .D(_03412_),
    .Q(\cpuregs[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27247_ (.CLK(clk),
    .D(_03413_),
    .Q(\cpuregs[3][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27248_ (.CLK(clk),
    .D(_03414_),
    .Q(\cpuregs[3][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27249_ (.CLK(clk),
    .D(_03415_),
    .Q(\cpuregs[3][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27250_ (.CLK(clk),
    .D(_03416_),
    .Q(\cpuregs[3][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27251_ (.CLK(clk),
    .D(_03417_),
    .Q(\cpuregs[3][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27252_ (.CLK(clk),
    .D(_03418_),
    .Q(\cpuregs[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27253_ (.CLK(clk),
    .D(_03419_),
    .Q(\cpuregs[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27254_ (.CLK(clk),
    .D(_03420_),
    .Q(\cpuregs[3][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27255_ (.CLK(clk),
    .D(_03421_),
    .Q(\cpuregs[3][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27256_ (.CLK(clk),
    .D(_03422_),
    .Q(\cpuregs[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27257_ (.CLK(clk),
    .D(_03423_),
    .Q(\cpuregs[3][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27258_ (.CLK(clk),
    .D(_03424_),
    .Q(\cpuregs[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27259_ (.CLK(clk),
    .D(_03425_),
    .Q(\cpuregs[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27260_ (.CLK(clk),
    .D(_03426_),
    .Q(\cpuregs[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27261_ (.CLK(clk),
    .D(_03427_),
    .Q(\cpuregs[3][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27262_ (.CLK(clk),
    .D(_03428_),
    .Q(\cpuregs[3][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27263_ (.CLK(clk),
    .D(_03429_),
    .Q(\cpuregs[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27264_ (.CLK(clk),
    .D(_03430_),
    .Q(\cpuregs[3][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27265_ (.CLK(clk),
    .D(_03431_),
    .Q(\cpuregs[3][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27266_ (.CLK(clk),
    .D(_03432_),
    .Q(\cpuregs[3][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27267_ (.CLK(clk),
    .D(_03433_),
    .Q(\cpuregs[3][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27268_ (.CLK(clk),
    .D(_03434_),
    .Q(\cpuregs[3][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27269_ (.CLK(clk),
    .D(_03435_),
    .Q(\cpuregs[3][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27270_ (.CLK(clk),
    .D(_03436_),
    .Q(\cpuregs[3][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27271_ (.CLK(clk),
    .D(_03437_),
    .Q(\cpuregs[3][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27272_ (.CLK(clk),
    .D(_03438_),
    .Q(\cpuregs[3][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27273_ (.CLK(clk),
    .D(_03439_),
    .Q(\cpuregs[11][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27274_ (.CLK(clk),
    .D(_03440_),
    .Q(\cpuregs[11][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27275_ (.CLK(clk),
    .D(_03441_),
    .Q(\cpuregs[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27276_ (.CLK(clk),
    .D(_03442_),
    .Q(\cpuregs[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27277_ (.CLK(clk),
    .D(_03443_),
    .Q(\cpuregs[11][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27278_ (.CLK(clk),
    .D(_03444_),
    .Q(\cpuregs[11][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27279_ (.CLK(clk),
    .D(_03445_),
    .Q(\cpuregs[11][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27280_ (.CLK(clk),
    .D(_03446_),
    .Q(\cpuregs[11][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27281_ (.CLK(clk),
    .D(_03447_),
    .Q(\cpuregs[11][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27282_ (.CLK(clk),
    .D(_03448_),
    .Q(\cpuregs[11][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27283_ (.CLK(clk),
    .D(_03449_),
    .Q(\cpuregs[11][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27284_ (.CLK(clk),
    .D(_03450_),
    .Q(\cpuregs[11][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27285_ (.CLK(clk),
    .D(_03451_),
    .Q(\cpuregs[11][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27286_ (.CLK(clk),
    .D(_03452_),
    .Q(\cpuregs[11][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27287_ (.CLK(clk),
    .D(_03453_),
    .Q(\cpuregs[11][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27288_ (.CLK(clk),
    .D(_03454_),
    .Q(\cpuregs[11][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27289_ (.CLK(clk),
    .D(_03455_),
    .Q(\cpuregs[11][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27290_ (.CLK(clk),
    .D(_03456_),
    .Q(\cpuregs[11][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27291_ (.CLK(clk),
    .D(_03457_),
    .Q(\cpuregs[11][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27292_ (.CLK(clk),
    .D(_03458_),
    .Q(\cpuregs[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27293_ (.CLK(clk),
    .D(_03459_),
    .Q(\cpuregs[11][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27294_ (.CLK(clk),
    .D(_03460_),
    .Q(\cpuregs[11][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27295_ (.CLK(clk),
    .D(_03461_),
    .Q(\cpuregs[11][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27296_ (.CLK(clk),
    .D(_03462_),
    .Q(\cpuregs[11][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27297_ (.CLK(clk),
    .D(_03463_),
    .Q(\cpuregs[11][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27298_ (.CLK(clk),
    .D(_03464_),
    .Q(\cpuregs[11][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27299_ (.CLK(clk),
    .D(_03465_),
    .Q(\cpuregs[11][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27300_ (.CLK(clk),
    .D(_03466_),
    .Q(\cpuregs[11][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27301_ (.CLK(clk),
    .D(_03467_),
    .Q(\cpuregs[11][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27302_ (.CLK(clk),
    .D(_03468_),
    .Q(\cpuregs[11][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27303_ (.CLK(clk),
    .D(_03469_),
    .Q(\cpuregs[11][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27304_ (.CLK(clk),
    .D(_03470_),
    .Q(\cpuregs[11][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27305_ (.CLK(clk),
    .D(_03471_),
    .Q(\cpuregs[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27306_ (.CLK(clk),
    .D(_03472_),
    .Q(\cpuregs[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27307_ (.CLK(clk),
    .D(_03473_),
    .Q(\cpuregs[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27308_ (.CLK(clk),
    .D(_03474_),
    .Q(\cpuregs[15][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27309_ (.CLK(clk),
    .D(_03475_),
    .Q(\cpuregs[15][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27310_ (.CLK(clk),
    .D(_03476_),
    .Q(\cpuregs[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27311_ (.CLK(clk),
    .D(_03477_),
    .Q(\cpuregs[15][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27312_ (.CLK(clk),
    .D(_03478_),
    .Q(\cpuregs[15][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27313_ (.CLK(clk),
    .D(_03479_),
    .Q(\cpuregs[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27314_ (.CLK(clk),
    .D(_03480_),
    .Q(\cpuregs[15][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27315_ (.CLK(clk),
    .D(_03481_),
    .Q(\cpuregs[15][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27316_ (.CLK(clk),
    .D(_03482_),
    .Q(\cpuregs[15][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27317_ (.CLK(clk),
    .D(_03483_),
    .Q(\cpuregs[15][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27318_ (.CLK(clk),
    .D(_03484_),
    .Q(\cpuregs[15][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27319_ (.CLK(clk),
    .D(_03485_),
    .Q(\cpuregs[15][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27320_ (.CLK(clk),
    .D(_03486_),
    .Q(\cpuregs[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27321_ (.CLK(clk),
    .D(_03487_),
    .Q(\cpuregs[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27322_ (.CLK(clk),
    .D(_03488_),
    .Q(\cpuregs[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27323_ (.CLK(clk),
    .D(_03489_),
    .Q(\cpuregs[15][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27324_ (.CLK(clk),
    .D(_03490_),
    .Q(\cpuregs[15][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27325_ (.CLK(clk),
    .D(_03491_),
    .Q(\cpuregs[15][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27326_ (.CLK(clk),
    .D(_03492_),
    .Q(\cpuregs[15][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27327_ (.CLK(clk),
    .D(_03493_),
    .Q(\cpuregs[15][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27328_ (.CLK(clk),
    .D(_03494_),
    .Q(\cpuregs[15][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27329_ (.CLK(clk),
    .D(_03495_),
    .Q(\cpuregs[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27330_ (.CLK(clk),
    .D(_03496_),
    .Q(\cpuregs[15][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27331_ (.CLK(clk),
    .D(_03497_),
    .Q(\cpuregs[15][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27332_ (.CLK(clk),
    .D(_03498_),
    .Q(\cpuregs[15][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27333_ (.CLK(clk),
    .D(_03499_),
    .Q(\cpuregs[15][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27334_ (.CLK(clk),
    .D(_03500_),
    .Q(\cpuregs[15][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27335_ (.CLK(clk),
    .D(_03501_),
    .Q(\cpuregs[15][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27336_ (.CLK(clk),
    .D(_03502_),
    .Q(\cpuregs[15][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27337_ (.CLK(clk),
    .D(_03503_),
    .Q(\latched_rd[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27338_ (.CLK(clk),
    .D(_03504_),
    .Q(\cpuregs[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27339_ (.CLK(clk),
    .D(_03505_),
    .Q(\cpuregs[7][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27340_ (.CLK(clk),
    .D(_03506_),
    .Q(\cpuregs[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27341_ (.CLK(clk),
    .D(_03507_),
    .Q(\cpuregs[7][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27342_ (.CLK(clk),
    .D(_03508_),
    .Q(\cpuregs[7][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27343_ (.CLK(clk),
    .D(_03509_),
    .Q(\cpuregs[7][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27344_ (.CLK(clk),
    .D(_03510_),
    .Q(\cpuregs[7][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27345_ (.CLK(clk),
    .D(_03511_),
    .Q(\cpuregs[7][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27346_ (.CLK(clk),
    .D(_03512_),
    .Q(\cpuregs[7][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27347_ (.CLK(clk),
    .D(_03513_),
    .Q(\cpuregs[7][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27348_ (.CLK(clk),
    .D(_03514_),
    .Q(\cpuregs[7][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27349_ (.CLK(clk),
    .D(_03515_),
    .Q(\cpuregs[7][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27350_ (.CLK(clk),
    .D(_03516_),
    .Q(\cpuregs[7][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27351_ (.CLK(clk),
    .D(_03517_),
    .Q(\cpuregs[7][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27352_ (.CLK(clk),
    .D(_03518_),
    .Q(\cpuregs[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27353_ (.CLK(clk),
    .D(_03519_),
    .Q(\cpuregs[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27354_ (.CLK(clk),
    .D(_03520_),
    .Q(\cpuregs[7][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27355_ (.CLK(clk),
    .D(_03521_),
    .Q(\cpuregs[7][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27356_ (.CLK(clk),
    .D(_03522_),
    .Q(\cpuregs[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27357_ (.CLK(clk),
    .D(_03523_),
    .Q(\cpuregs[7][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27358_ (.CLK(clk),
    .D(_03524_),
    .Q(\cpuregs[7][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27359_ (.CLK(clk),
    .D(_03525_),
    .Q(\cpuregs[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27360_ (.CLK(clk),
    .D(_03526_),
    .Q(\cpuregs[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27361_ (.CLK(clk),
    .D(_03527_),
    .Q(\cpuregs[7][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27362_ (.CLK(clk),
    .D(_03528_),
    .Q(\cpuregs[7][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27363_ (.CLK(clk),
    .D(_03529_),
    .Q(\cpuregs[7][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27364_ (.CLK(clk),
    .D(_03530_),
    .Q(\cpuregs[7][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27365_ (.CLK(clk),
    .D(_03531_),
    .Q(\cpuregs[7][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27366_ (.CLK(clk),
    .D(_03532_),
    .Q(\cpuregs[7][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27367_ (.CLK(clk),
    .D(_03533_),
    .Q(\cpuregs[7][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27368_ (.CLK(clk),
    .D(_03534_),
    .Q(\cpuregs[7][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27369_ (.CLK(clk),
    .D(_03535_),
    .Q(\cpuregs[7][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27370_ (.CLK(clk),
    .D(_03536_),
    .Q(mem_wdata[0]));
 sky130_fd_sc_hd__dfxtp_2 _27371_ (.CLK(clk),
    .D(_03537_),
    .Q(mem_wdata[1]));
 sky130_fd_sc_hd__dfxtp_2 _27372_ (.CLK(clk),
    .D(_03538_),
    .Q(mem_wdata[2]));
 sky130_fd_sc_hd__dfxtp_2 _27373_ (.CLK(clk),
    .D(_03539_),
    .Q(mem_wdata[3]));
 sky130_fd_sc_hd__dfxtp_2 _27374_ (.CLK(clk),
    .D(_03540_),
    .Q(mem_wdata[4]));
 sky130_fd_sc_hd__dfxtp_2 _27375_ (.CLK(clk),
    .D(_03541_),
    .Q(mem_wdata[5]));
 sky130_fd_sc_hd__dfxtp_2 _27376_ (.CLK(clk),
    .D(_03542_),
    .Q(mem_wdata[6]));
 sky130_fd_sc_hd__dfxtp_2 _27377_ (.CLK(clk),
    .D(_03543_),
    .Q(mem_wdata[7]));
 sky130_fd_sc_hd__dfxtp_2 _27378_ (.CLK(clk),
    .D(_03544_),
    .Q(mem_wdata[8]));
 sky130_fd_sc_hd__dfxtp_2 _27379_ (.CLK(clk),
    .D(_03545_),
    .Q(mem_wdata[9]));
 sky130_fd_sc_hd__dfxtp_2 _27380_ (.CLK(clk),
    .D(_03546_),
    .Q(mem_wdata[10]));
 sky130_fd_sc_hd__dfxtp_2 _27381_ (.CLK(clk),
    .D(_03547_),
    .Q(mem_wdata[11]));
 sky130_fd_sc_hd__dfxtp_2 _27382_ (.CLK(clk),
    .D(_03548_),
    .Q(mem_wdata[12]));
 sky130_fd_sc_hd__dfxtp_2 _27383_ (.CLK(clk),
    .D(_03549_),
    .Q(mem_wdata[13]));
 sky130_fd_sc_hd__dfxtp_2 _27384_ (.CLK(clk),
    .D(_03550_),
    .Q(mem_wdata[14]));
 sky130_fd_sc_hd__dfxtp_2 _27385_ (.CLK(clk),
    .D(_03551_),
    .Q(mem_wdata[15]));
 sky130_fd_sc_hd__dfxtp_2 _27386_ (.CLK(clk),
    .D(_03552_),
    .Q(mem_wdata[16]));
 sky130_fd_sc_hd__dfxtp_2 _27387_ (.CLK(clk),
    .D(_03553_),
    .Q(mem_wdata[17]));
 sky130_fd_sc_hd__dfxtp_2 _27388_ (.CLK(clk),
    .D(_03554_),
    .Q(mem_wdata[18]));
 sky130_fd_sc_hd__dfxtp_2 _27389_ (.CLK(clk),
    .D(_03555_),
    .Q(mem_wdata[19]));
 sky130_fd_sc_hd__dfxtp_2 _27390_ (.CLK(clk),
    .D(_03556_),
    .Q(mem_wdata[20]));
 sky130_fd_sc_hd__dfxtp_2 _27391_ (.CLK(clk),
    .D(_03557_),
    .Q(mem_wdata[21]));
 sky130_fd_sc_hd__dfxtp_2 _27392_ (.CLK(clk),
    .D(_03558_),
    .Q(mem_wdata[22]));
 sky130_fd_sc_hd__dfxtp_2 _27393_ (.CLK(clk),
    .D(_03559_),
    .Q(mem_wdata[23]));
 sky130_fd_sc_hd__dfxtp_2 _27394_ (.CLK(clk),
    .D(_03560_),
    .Q(mem_wdata[24]));
 sky130_fd_sc_hd__dfxtp_2 _27395_ (.CLK(clk),
    .D(_03561_),
    .Q(mem_wdata[25]));
 sky130_fd_sc_hd__dfxtp_2 _27396_ (.CLK(clk),
    .D(_03562_),
    .Q(mem_wdata[26]));
 sky130_fd_sc_hd__dfxtp_2 _27397_ (.CLK(clk),
    .D(_03563_),
    .Q(mem_wdata[27]));
 sky130_fd_sc_hd__dfxtp_2 _27398_ (.CLK(clk),
    .D(_03564_),
    .Q(mem_wdata[28]));
 sky130_fd_sc_hd__dfxtp_2 _27399_ (.CLK(clk),
    .D(_03565_),
    .Q(mem_wdata[29]));
 sky130_fd_sc_hd__dfxtp_2 _27400_ (.CLK(clk),
    .D(_03566_),
    .Q(mem_wdata[30]));
 sky130_fd_sc_hd__dfxtp_2 _27401_ (.CLK(clk),
    .D(_03567_),
    .Q(mem_wdata[31]));
 sky130_fd_sc_hd__dfxtp_2 _27402_ (.CLK(clk),
    .D(_03568_),
    .Q(\cpuregs[19][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27403_ (.CLK(clk),
    .D(_03569_),
    .Q(\cpuregs[19][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27404_ (.CLK(clk),
    .D(_03570_),
    .Q(\cpuregs[19][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27405_ (.CLK(clk),
    .D(_03571_),
    .Q(\cpuregs[19][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27406_ (.CLK(clk),
    .D(_03572_),
    .Q(\cpuregs[19][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27407_ (.CLK(clk),
    .D(_03573_),
    .Q(\cpuregs[19][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27408_ (.CLK(clk),
    .D(_03574_),
    .Q(\cpuregs[19][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27409_ (.CLK(clk),
    .D(_03575_),
    .Q(\cpuregs[19][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27410_ (.CLK(clk),
    .D(_03576_),
    .Q(\cpuregs[19][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27411_ (.CLK(clk),
    .D(_03577_),
    .Q(\cpuregs[19][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27412_ (.CLK(clk),
    .D(_03578_),
    .Q(\cpuregs[19][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27413_ (.CLK(clk),
    .D(_03579_),
    .Q(\cpuregs[19][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27414_ (.CLK(clk),
    .D(_03580_),
    .Q(\cpuregs[19][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27415_ (.CLK(clk),
    .D(_03581_),
    .Q(\cpuregs[19][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27416_ (.CLK(clk),
    .D(_03582_),
    .Q(\cpuregs[19][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27417_ (.CLK(clk),
    .D(_03583_),
    .Q(\cpuregs[19][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27418_ (.CLK(clk),
    .D(_03584_),
    .Q(\cpuregs[19][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27419_ (.CLK(clk),
    .D(_03585_),
    .Q(\cpuregs[19][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27420_ (.CLK(clk),
    .D(_03586_),
    .Q(\cpuregs[19][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27421_ (.CLK(clk),
    .D(_03587_),
    .Q(\cpuregs[19][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27422_ (.CLK(clk),
    .D(_03588_),
    .Q(\cpuregs[19][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27423_ (.CLK(clk),
    .D(_03589_),
    .Q(\cpuregs[19][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27424_ (.CLK(clk),
    .D(_03590_),
    .Q(\cpuregs[19][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27425_ (.CLK(clk),
    .D(_03591_),
    .Q(\cpuregs[19][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27426_ (.CLK(clk),
    .D(_03592_),
    .Q(\cpuregs[19][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27427_ (.CLK(clk),
    .D(_03593_),
    .Q(\cpuregs[19][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27428_ (.CLK(clk),
    .D(_03594_),
    .Q(\cpuregs[19][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27429_ (.CLK(clk),
    .D(_03595_),
    .Q(\cpuregs[19][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27430_ (.CLK(clk),
    .D(_03596_),
    .Q(\cpuregs[19][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27431_ (.CLK(clk),
    .D(_03597_),
    .Q(\cpuregs[19][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27432_ (.CLK(clk),
    .D(_03598_),
    .Q(\cpuregs[19][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27433_ (.CLK(clk),
    .D(_03599_),
    .Q(\cpuregs[19][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27434_ (.CLK(clk),
    .D(_03600_),
    .Q(\cpuregs[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27435_ (.CLK(clk),
    .D(_03601_),
    .Q(\cpuregs[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27436_ (.CLK(clk),
    .D(_03602_),
    .Q(\cpuregs[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27437_ (.CLK(clk),
    .D(_03603_),
    .Q(\cpuregs[4][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27438_ (.CLK(clk),
    .D(_03604_),
    .Q(\cpuregs[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27439_ (.CLK(clk),
    .D(_03605_),
    .Q(\cpuregs[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27440_ (.CLK(clk),
    .D(_03606_),
    .Q(\cpuregs[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27441_ (.CLK(clk),
    .D(_03607_),
    .Q(\cpuregs[4][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27442_ (.CLK(clk),
    .D(_03608_),
    .Q(\cpuregs[4][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27443_ (.CLK(clk),
    .D(_03609_),
    .Q(\cpuregs[4][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27444_ (.CLK(clk),
    .D(_03610_),
    .Q(\cpuregs[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27445_ (.CLK(clk),
    .D(_03611_),
    .Q(\cpuregs[4][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27446_ (.CLK(clk),
    .D(_03612_),
    .Q(\cpuregs[4][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27447_ (.CLK(clk),
    .D(_03613_),
    .Q(\cpuregs[4][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27448_ (.CLK(clk),
    .D(_03614_),
    .Q(\cpuregs[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27449_ (.CLK(clk),
    .D(_03615_),
    .Q(\cpuregs[4][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27450_ (.CLK(clk),
    .D(_03616_),
    .Q(\cpuregs[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27451_ (.CLK(clk),
    .D(_03617_),
    .Q(\cpuregs[4][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27452_ (.CLK(clk),
    .D(_03618_),
    .Q(\cpuregs[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27453_ (.CLK(clk),
    .D(_03619_),
    .Q(\cpuregs[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27454_ (.CLK(clk),
    .D(_03620_),
    .Q(\cpuregs[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27455_ (.CLK(clk),
    .D(_03621_),
    .Q(\cpuregs[4][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27456_ (.CLK(clk),
    .D(_03622_),
    .Q(\cpuregs[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27457_ (.CLK(clk),
    .D(_03623_),
    .Q(\cpuregs[4][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27458_ (.CLK(clk),
    .D(_03624_),
    .Q(\cpuregs[4][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27459_ (.CLK(clk),
    .D(_03625_),
    .Q(\cpuregs[4][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27460_ (.CLK(clk),
    .D(_03626_),
    .Q(\cpuregs[4][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27461_ (.CLK(clk),
    .D(_03627_),
    .Q(\cpuregs[4][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27462_ (.CLK(clk),
    .D(_03628_),
    .Q(\cpuregs[4][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27463_ (.CLK(clk),
    .D(_03629_),
    .Q(\cpuregs[4][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27464_ (.CLK(clk),
    .D(_03630_),
    .Q(\cpuregs[4][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27465_ (.CLK(clk),
    .D(_03631_),
    .Q(\cpuregs[4][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27466_ (.CLK(clk),
    .D(_03632_),
    .Q(mem_la_wdata[0]));
 sky130_fd_sc_hd__dfxtp_2 _27467_ (.CLK(clk),
    .D(_03633_),
    .Q(mem_la_wdata[1]));
 sky130_fd_sc_hd__dfxtp_2 _27468_ (.CLK(clk),
    .D(_03634_),
    .Q(mem_la_wdata[2]));
 sky130_fd_sc_hd__dfxtp_2 _27469_ (.CLK(clk),
    .D(_03635_),
    .Q(mem_la_wdata[3]));
 sky130_fd_sc_hd__dfxtp_2 _27470_ (.CLK(clk),
    .D(_03636_),
    .Q(mem_la_wdata[4]));
 sky130_fd_sc_hd__dfxtp_2 _27471_ (.CLK(clk),
    .D(_03637_),
    .Q(mem_la_wdata[5]));
 sky130_fd_sc_hd__dfxtp_2 _27472_ (.CLK(clk),
    .D(_03638_),
    .Q(mem_la_wdata[6]));
 sky130_fd_sc_hd__dfxtp_2 _27473_ (.CLK(clk),
    .D(_03639_),
    .Q(mem_la_wdata[7]));
 sky130_fd_sc_hd__dfxtp_2 _27474_ (.CLK(clk),
    .D(_03640_),
    .Q(pcpi_rs2[8]));
 sky130_fd_sc_hd__dfxtp_2 _27475_ (.CLK(clk),
    .D(_03641_),
    .Q(pcpi_rs2[9]));
 sky130_fd_sc_hd__dfxtp_2 _27476_ (.CLK(clk),
    .D(_03642_),
    .Q(pcpi_rs2[10]));
 sky130_fd_sc_hd__dfxtp_2 _27477_ (.CLK(clk),
    .D(_03643_),
    .Q(pcpi_rs2[11]));
 sky130_fd_sc_hd__dfxtp_2 _27478_ (.CLK(clk),
    .D(_03644_),
    .Q(pcpi_rs2[12]));
 sky130_fd_sc_hd__dfxtp_2 _27479_ (.CLK(clk),
    .D(_03645_),
    .Q(pcpi_rs2[13]));
 sky130_fd_sc_hd__dfxtp_2 _27480_ (.CLK(clk),
    .D(_03646_),
    .Q(pcpi_rs2[14]));
 sky130_fd_sc_hd__dfxtp_2 _27481_ (.CLK(clk),
    .D(_03647_),
    .Q(pcpi_rs2[15]));
 sky130_fd_sc_hd__dfxtp_2 _27482_ (.CLK(clk),
    .D(_03648_),
    .Q(pcpi_rs2[16]));
 sky130_fd_sc_hd__dfxtp_2 _27483_ (.CLK(clk),
    .D(_03649_),
    .Q(pcpi_rs2[17]));
 sky130_fd_sc_hd__dfxtp_2 _27484_ (.CLK(clk),
    .D(_03650_),
    .Q(pcpi_rs2[18]));
 sky130_fd_sc_hd__dfxtp_2 _27485_ (.CLK(clk),
    .D(_03651_),
    .Q(pcpi_rs2[19]));
 sky130_fd_sc_hd__dfxtp_2 _27486_ (.CLK(clk),
    .D(_03652_),
    .Q(pcpi_rs2[20]));
 sky130_fd_sc_hd__dfxtp_2 _27487_ (.CLK(clk),
    .D(_03653_),
    .Q(pcpi_rs2[21]));
 sky130_fd_sc_hd__dfxtp_2 _27488_ (.CLK(clk),
    .D(_03654_),
    .Q(pcpi_rs2[22]));
 sky130_fd_sc_hd__dfxtp_2 _27489_ (.CLK(clk),
    .D(_03655_),
    .Q(pcpi_rs2[23]));
 sky130_fd_sc_hd__dfxtp_2 _27490_ (.CLK(clk),
    .D(_03656_),
    .Q(pcpi_rs2[24]));
 sky130_fd_sc_hd__dfxtp_2 _27491_ (.CLK(clk),
    .D(_03657_),
    .Q(pcpi_rs2[25]));
 sky130_fd_sc_hd__dfxtp_2 _27492_ (.CLK(clk),
    .D(_03658_),
    .Q(pcpi_rs2[26]));
 sky130_fd_sc_hd__dfxtp_2 _27493_ (.CLK(clk),
    .D(_03659_),
    .Q(pcpi_rs2[27]));
 sky130_fd_sc_hd__dfxtp_2 _27494_ (.CLK(clk),
    .D(_03660_),
    .Q(pcpi_rs2[28]));
 sky130_fd_sc_hd__dfxtp_2 _27495_ (.CLK(clk),
    .D(_03661_),
    .Q(pcpi_rs2[29]));
 sky130_fd_sc_hd__dfxtp_2 _27496_ (.CLK(clk),
    .D(_03662_),
    .Q(pcpi_rs2[30]));
 sky130_fd_sc_hd__dfxtp_2 _27497_ (.CLK(clk),
    .D(_03663_),
    .Q(pcpi_rs2[31]));
 sky130_fd_sc_hd__dfxtp_2 _27498_ (.CLK(clk),
    .D(_03664_),
    .Q(\cpuregs[9][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27499_ (.CLK(clk),
    .D(_03665_),
    .Q(\cpuregs[9][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27500_ (.CLK(clk),
    .D(_03666_),
    .Q(\cpuregs[9][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27501_ (.CLK(clk),
    .D(_03667_),
    .Q(\cpuregs[9][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27502_ (.CLK(clk),
    .D(_03668_),
    .Q(\cpuregs[9][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27503_ (.CLK(clk),
    .D(_03669_),
    .Q(\cpuregs[9][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27504_ (.CLK(clk),
    .D(_03670_),
    .Q(\cpuregs[9][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27505_ (.CLK(clk),
    .D(_03671_),
    .Q(\cpuregs[9][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27506_ (.CLK(clk),
    .D(_03672_),
    .Q(\cpuregs[9][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27507_ (.CLK(clk),
    .D(_03673_),
    .Q(\cpuregs[9][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27508_ (.CLK(clk),
    .D(_03674_),
    .Q(\cpuregs[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27509_ (.CLK(clk),
    .D(_03675_),
    .Q(\cpuregs[9][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27510_ (.CLK(clk),
    .D(_03676_),
    .Q(\cpuregs[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27511_ (.CLK(clk),
    .D(_03677_),
    .Q(\cpuregs[9][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27512_ (.CLK(clk),
    .D(_03678_),
    .Q(\cpuregs[9][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27513_ (.CLK(clk),
    .D(_03679_),
    .Q(\cpuregs[9][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27514_ (.CLK(clk),
    .D(_03680_),
    .Q(\cpuregs[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27515_ (.CLK(clk),
    .D(_03681_),
    .Q(\cpuregs[9][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27516_ (.CLK(clk),
    .D(_03682_),
    .Q(\cpuregs[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27517_ (.CLK(clk),
    .D(_03683_),
    .Q(\cpuregs[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27518_ (.CLK(clk),
    .D(_03684_),
    .Q(\cpuregs[9][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27519_ (.CLK(clk),
    .D(_03685_),
    .Q(\cpuregs[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27520_ (.CLK(clk),
    .D(_03686_),
    .Q(\cpuregs[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27521_ (.CLK(clk),
    .D(_03687_),
    .Q(\cpuregs[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27522_ (.CLK(clk),
    .D(_03688_),
    .Q(\cpuregs[9][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27523_ (.CLK(clk),
    .D(_03689_),
    .Q(\cpuregs[9][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27524_ (.CLK(clk),
    .D(_03690_),
    .Q(\cpuregs[9][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27525_ (.CLK(clk),
    .D(_03691_),
    .Q(\cpuregs[9][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27526_ (.CLK(clk),
    .D(_03692_),
    .Q(\cpuregs[9][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27527_ (.CLK(clk),
    .D(_03693_),
    .Q(\cpuregs[9][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27528_ (.CLK(clk),
    .D(_03694_),
    .Q(\cpuregs[9][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27529_ (.CLK(clk),
    .D(_03695_),
    .Q(\cpuregs[9][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27530_ (.CLK(clk),
    .D(_03696_),
    .Q(\cpuregs[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _27531_ (.CLK(clk),
    .D(_03697_),
    .Q(\cpuregs[6][1] ));
 sky130_fd_sc_hd__dfxtp_2 _27532_ (.CLK(clk),
    .D(_03698_),
    .Q(\cpuregs[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _27533_ (.CLK(clk),
    .D(_03699_),
    .Q(\cpuregs[6][3] ));
 sky130_fd_sc_hd__dfxtp_2 _27534_ (.CLK(clk),
    .D(_03700_),
    .Q(\cpuregs[6][4] ));
 sky130_fd_sc_hd__dfxtp_2 _27535_ (.CLK(clk),
    .D(_03701_),
    .Q(\cpuregs[6][5] ));
 sky130_fd_sc_hd__dfxtp_2 _27536_ (.CLK(clk),
    .D(_03702_),
    .Q(\cpuregs[6][6] ));
 sky130_fd_sc_hd__dfxtp_2 _27537_ (.CLK(clk),
    .D(_03703_),
    .Q(\cpuregs[6][7] ));
 sky130_fd_sc_hd__dfxtp_2 _27538_ (.CLK(clk),
    .D(_03704_),
    .Q(\cpuregs[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _27539_ (.CLK(clk),
    .D(_03705_),
    .Q(\cpuregs[6][9] ));
 sky130_fd_sc_hd__dfxtp_2 _27540_ (.CLK(clk),
    .D(_03706_),
    .Q(\cpuregs[6][10] ));
 sky130_fd_sc_hd__dfxtp_2 _27541_ (.CLK(clk),
    .D(_03707_),
    .Q(\cpuregs[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _27542_ (.CLK(clk),
    .D(_03708_),
    .Q(\cpuregs[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _27543_ (.CLK(clk),
    .D(_03709_),
    .Q(\cpuregs[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _27544_ (.CLK(clk),
    .D(_03710_),
    .Q(\cpuregs[6][14] ));
 sky130_fd_sc_hd__dfxtp_2 _27545_ (.CLK(clk),
    .D(_03711_),
    .Q(\cpuregs[6][15] ));
 sky130_fd_sc_hd__dfxtp_2 _27546_ (.CLK(clk),
    .D(_03712_),
    .Q(\cpuregs[6][16] ));
 sky130_fd_sc_hd__dfxtp_2 _27547_ (.CLK(clk),
    .D(_03713_),
    .Q(\cpuregs[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _27548_ (.CLK(clk),
    .D(_03714_),
    .Q(\cpuregs[6][18] ));
 sky130_fd_sc_hd__dfxtp_2 _27549_ (.CLK(clk),
    .D(_03715_),
    .Q(\cpuregs[6][19] ));
 sky130_fd_sc_hd__dfxtp_2 _27550_ (.CLK(clk),
    .D(_03716_),
    .Q(\cpuregs[6][20] ));
 sky130_fd_sc_hd__dfxtp_2 _27551_ (.CLK(clk),
    .D(_03717_),
    .Q(\cpuregs[6][21] ));
 sky130_fd_sc_hd__dfxtp_2 _27552_ (.CLK(clk),
    .D(_03718_),
    .Q(\cpuregs[6][22] ));
 sky130_fd_sc_hd__dfxtp_2 _27553_ (.CLK(clk),
    .D(_03719_),
    .Q(\cpuregs[6][23] ));
 sky130_fd_sc_hd__dfxtp_2 _27554_ (.CLK(clk),
    .D(_03720_),
    .Q(\cpuregs[6][24] ));
 sky130_fd_sc_hd__dfxtp_2 _27555_ (.CLK(clk),
    .D(_03721_),
    .Q(\cpuregs[6][25] ));
 sky130_fd_sc_hd__dfxtp_2 _27556_ (.CLK(clk),
    .D(_03722_),
    .Q(\cpuregs[6][26] ));
 sky130_fd_sc_hd__dfxtp_2 _27557_ (.CLK(clk),
    .D(_03723_),
    .Q(\cpuregs[6][27] ));
 sky130_fd_sc_hd__dfxtp_2 _27558_ (.CLK(clk),
    .D(_03724_),
    .Q(\cpuregs[6][28] ));
 sky130_fd_sc_hd__dfxtp_2 _27559_ (.CLK(clk),
    .D(_03725_),
    .Q(\cpuregs[6][29] ));
 sky130_fd_sc_hd__dfxtp_2 _27560_ (.CLK(clk),
    .D(_03726_),
    .Q(\cpuregs[6][30] ));
 sky130_fd_sc_hd__dfxtp_2 _27561_ (.CLK(clk),
    .D(_03727_),
    .Q(\cpuregs[6][31] ));
 sky130_fd_sc_hd__dfxtp_2 _27562_ (.CLK(clk),
    .D(_03728_),
    .Q(\pcpi_mul.active[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27563_ (.CLK(clk),
    .D(_03729_),
    .Q(\pcpi_mul.active[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27564_ (.CLK(clk),
    .D(_03730_),
    .Q(trap));
 sky130_fd_sc_hd__dfxtp_2 _27565_ (.CLK(clk),
    .D(_03731_),
    .Q(\count_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27566_ (.CLK(clk),
    .D(_03732_),
    .Q(\count_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27567_ (.CLK(clk),
    .D(_03733_),
    .Q(\count_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27568_ (.CLK(clk),
    .D(_03734_),
    .Q(\count_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27569_ (.CLK(clk),
    .D(_03735_),
    .Q(\count_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27570_ (.CLK(clk),
    .D(_03736_),
    .Q(\count_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27571_ (.CLK(clk),
    .D(_03737_),
    .Q(\count_cycle[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27572_ (.CLK(clk),
    .D(_03738_),
    .Q(\count_cycle[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27573_ (.CLK(clk),
    .D(_03739_),
    .Q(\count_cycle[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27574_ (.CLK(clk),
    .D(_03740_),
    .Q(\count_cycle[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27575_ (.CLK(clk),
    .D(_03741_),
    .Q(\count_cycle[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27576_ (.CLK(clk),
    .D(_03742_),
    .Q(\count_cycle[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27577_ (.CLK(clk),
    .D(_03743_),
    .Q(\count_cycle[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27578_ (.CLK(clk),
    .D(_03744_),
    .Q(\count_cycle[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27579_ (.CLK(clk),
    .D(_03745_),
    .Q(\count_cycle[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27580_ (.CLK(clk),
    .D(_03746_),
    .Q(\count_cycle[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27581_ (.CLK(clk),
    .D(_03747_),
    .Q(\count_cycle[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27582_ (.CLK(clk),
    .D(_03748_),
    .Q(\count_cycle[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27583_ (.CLK(clk),
    .D(_03749_),
    .Q(\count_cycle[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27584_ (.CLK(clk),
    .D(_03750_),
    .Q(\count_cycle[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27585_ (.CLK(clk),
    .D(_03751_),
    .Q(\count_cycle[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27586_ (.CLK(clk),
    .D(_03752_),
    .Q(\count_cycle[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27587_ (.CLK(clk),
    .D(_03753_),
    .Q(\count_cycle[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27588_ (.CLK(clk),
    .D(_03754_),
    .Q(\count_cycle[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27589_ (.CLK(clk),
    .D(_03755_),
    .Q(\count_cycle[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27590_ (.CLK(clk),
    .D(_03756_),
    .Q(\count_cycle[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27591_ (.CLK(clk),
    .D(_03757_),
    .Q(\count_cycle[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27592_ (.CLK(clk),
    .D(_03758_),
    .Q(\count_cycle[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27593_ (.CLK(clk),
    .D(_03759_),
    .Q(\count_cycle[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27594_ (.CLK(clk),
    .D(_03760_),
    .Q(\count_cycle[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27595_ (.CLK(clk),
    .D(_03761_),
    .Q(\count_cycle[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27596_ (.CLK(clk),
    .D(_03762_),
    .Q(\count_cycle[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27597_ (.CLK(clk),
    .D(_03763_),
    .Q(\count_cycle[32] ));
 sky130_fd_sc_hd__dfxtp_2 _27598_ (.CLK(clk),
    .D(_03764_),
    .Q(\count_cycle[33] ));
 sky130_fd_sc_hd__dfxtp_2 _27599_ (.CLK(clk),
    .D(_03765_),
    .Q(\count_cycle[34] ));
 sky130_fd_sc_hd__dfxtp_2 _27600_ (.CLK(clk),
    .D(_03766_),
    .Q(\count_cycle[35] ));
 sky130_fd_sc_hd__dfxtp_2 _27601_ (.CLK(clk),
    .D(_03767_),
    .Q(\count_cycle[36] ));
 sky130_fd_sc_hd__dfxtp_2 _27602_ (.CLK(clk),
    .D(_03768_),
    .Q(\count_cycle[37] ));
 sky130_fd_sc_hd__dfxtp_2 _27603_ (.CLK(clk),
    .D(_03769_),
    .Q(\count_cycle[38] ));
 sky130_fd_sc_hd__dfxtp_2 _27604_ (.CLK(clk),
    .D(_03770_),
    .Q(\count_cycle[39] ));
 sky130_fd_sc_hd__dfxtp_2 _27605_ (.CLK(clk),
    .D(_03771_),
    .Q(\count_cycle[40] ));
 sky130_fd_sc_hd__dfxtp_2 _27606_ (.CLK(clk),
    .D(_03772_),
    .Q(\count_cycle[41] ));
 sky130_fd_sc_hd__dfxtp_2 _27607_ (.CLK(clk),
    .D(_03773_),
    .Q(\count_cycle[42] ));
 sky130_fd_sc_hd__dfxtp_2 _27608_ (.CLK(clk),
    .D(_03774_),
    .Q(\count_cycle[43] ));
 sky130_fd_sc_hd__dfxtp_2 _27609_ (.CLK(clk),
    .D(_03775_),
    .Q(\count_cycle[44] ));
 sky130_fd_sc_hd__dfxtp_2 _27610_ (.CLK(clk),
    .D(_03776_),
    .Q(\count_cycle[45] ));
 sky130_fd_sc_hd__dfxtp_2 _27611_ (.CLK(clk),
    .D(_03777_),
    .Q(\count_cycle[46] ));
 sky130_fd_sc_hd__dfxtp_2 _27612_ (.CLK(clk),
    .D(_03778_),
    .Q(\count_cycle[47] ));
 sky130_fd_sc_hd__dfxtp_2 _27613_ (.CLK(clk),
    .D(_03779_),
    .Q(\count_cycle[48] ));
 sky130_fd_sc_hd__dfxtp_2 _27614_ (.CLK(clk),
    .D(_03780_),
    .Q(\count_cycle[49] ));
 sky130_fd_sc_hd__dfxtp_2 _27615_ (.CLK(clk),
    .D(_03781_),
    .Q(\count_cycle[50] ));
 sky130_fd_sc_hd__dfxtp_2 _27616_ (.CLK(clk),
    .D(_03782_),
    .Q(\count_cycle[51] ));
 sky130_fd_sc_hd__dfxtp_2 _27617_ (.CLK(clk),
    .D(_03783_),
    .Q(\count_cycle[52] ));
 sky130_fd_sc_hd__dfxtp_2 _27618_ (.CLK(clk),
    .D(_03784_),
    .Q(\count_cycle[53] ));
 sky130_fd_sc_hd__dfxtp_2 _27619_ (.CLK(clk),
    .D(_03785_),
    .Q(\count_cycle[54] ));
 sky130_fd_sc_hd__dfxtp_2 _27620_ (.CLK(clk),
    .D(_03786_),
    .Q(\count_cycle[55] ));
 sky130_fd_sc_hd__dfxtp_2 _27621_ (.CLK(clk),
    .D(_03787_),
    .Q(\count_cycle[56] ));
 sky130_fd_sc_hd__dfxtp_2 _27622_ (.CLK(clk),
    .D(_03788_),
    .Q(\count_cycle[57] ));
 sky130_fd_sc_hd__dfxtp_2 _27623_ (.CLK(clk),
    .D(_03789_),
    .Q(\count_cycle[58] ));
 sky130_fd_sc_hd__dfxtp_2 _27624_ (.CLK(clk),
    .D(_03790_),
    .Q(\count_cycle[59] ));
 sky130_fd_sc_hd__dfxtp_2 _27625_ (.CLK(clk),
    .D(_03791_),
    .Q(\count_cycle[60] ));
 sky130_fd_sc_hd__dfxtp_2 _27626_ (.CLK(clk),
    .D(_03792_),
    .Q(\count_cycle[61] ));
 sky130_fd_sc_hd__dfxtp_2 _27627_ (.CLK(clk),
    .D(_03793_),
    .Q(\count_cycle[62] ));
 sky130_fd_sc_hd__dfxtp_2 _27628_ (.CLK(clk),
    .D(_03794_),
    .Q(\count_cycle[63] ));
 sky130_fd_sc_hd__dfxtp_2 _27629_ (.CLK(clk),
    .D(_03795_),
    .Q(\timer[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27630_ (.CLK(clk),
    .D(_03796_),
    .Q(\timer[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27631_ (.CLK(clk),
    .D(_03797_),
    .Q(\timer[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27632_ (.CLK(clk),
    .D(_03798_),
    .Q(\timer[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27633_ (.CLK(clk),
    .D(_03799_),
    .Q(\timer[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27634_ (.CLK(clk),
    .D(_03800_),
    .Q(\timer[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27635_ (.CLK(clk),
    .D(_03801_),
    .Q(\timer[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27636_ (.CLK(clk),
    .D(_03802_),
    .Q(\timer[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27637_ (.CLK(clk),
    .D(_03803_),
    .Q(\timer[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27638_ (.CLK(clk),
    .D(_03804_),
    .Q(\timer[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27639_ (.CLK(clk),
    .D(_03805_),
    .Q(\timer[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27640_ (.CLK(clk),
    .D(_03806_),
    .Q(\timer[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27641_ (.CLK(clk),
    .D(_03807_),
    .Q(\timer[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27642_ (.CLK(clk),
    .D(_03808_),
    .Q(\timer[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27643_ (.CLK(clk),
    .D(_03809_),
    .Q(\timer[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27644_ (.CLK(clk),
    .D(_03810_),
    .Q(\timer[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27645_ (.CLK(clk),
    .D(_03811_),
    .Q(\timer[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27646_ (.CLK(clk),
    .D(_03812_),
    .Q(\timer[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27647_ (.CLK(clk),
    .D(_03813_),
    .Q(\timer[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27648_ (.CLK(clk),
    .D(_03814_),
    .Q(\timer[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27649_ (.CLK(clk),
    .D(_03815_),
    .Q(\timer[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27650_ (.CLK(clk),
    .D(_03816_),
    .Q(\timer[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27651_ (.CLK(clk),
    .D(_03817_),
    .Q(\timer[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27652_ (.CLK(clk),
    .D(_03818_),
    .Q(\timer[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27653_ (.CLK(clk),
    .D(_03819_),
    .Q(\timer[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27654_ (.CLK(clk),
    .D(_03820_),
    .Q(\timer[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27655_ (.CLK(clk),
    .D(_03821_),
    .Q(\timer[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27656_ (.CLK(clk),
    .D(_03822_),
    .Q(\timer[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27657_ (.CLK(clk),
    .D(_03823_),
    .Q(\timer[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27658_ (.CLK(clk),
    .D(_03824_),
    .Q(\timer[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27659_ (.CLK(clk),
    .D(_03825_),
    .Q(\timer[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27660_ (.CLK(clk),
    .D(_03826_),
    .Q(\timer[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27661_ (.CLK(clk),
    .D(_03827_),
    .Q(pcpi_timeout));
 sky130_fd_sc_hd__dfxtp_2 _27662_ (.CLK(clk),
    .D(_03828_),
    .Q(decoder_pseudo_trigger));
 sky130_fd_sc_hd__dfxtp_2 _27663_ (.CLK(clk),
    .D(_03829_),
    .Q(is_compare));
 sky130_fd_sc_hd__dfxtp_2 _27664_ (.CLK(clk),
    .D(_03830_),
    .Q(do_waitirq));
 sky130_fd_sc_hd__dfxtp_2 _27665_ (.CLK(clk),
    .D(_03831_),
    .Q(mem_valid));
 sky130_fd_sc_hd__dfxtp_2 _27666_ (.CLK(clk),
    .D(_03832_),
    .Q(pcpi_valid));
 sky130_fd_sc_hd__dfxtp_2 _27667_ (.CLK(clk),
    .D(_03833_),
    .Q(eoi[0]));
 sky130_fd_sc_hd__dfxtp_2 _27668_ (.CLK(clk),
    .D(_03834_),
    .Q(eoi[1]));
 sky130_fd_sc_hd__dfxtp_2 _27669_ (.CLK(clk),
    .D(_03835_),
    .Q(eoi[2]));
 sky130_fd_sc_hd__dfxtp_2 _27670_ (.CLK(clk),
    .D(_03836_),
    .Q(eoi[3]));
 sky130_fd_sc_hd__dfxtp_2 _27671_ (.CLK(clk),
    .D(_03837_),
    .Q(eoi[4]));
 sky130_fd_sc_hd__dfxtp_2 _27672_ (.CLK(clk),
    .D(_03838_),
    .Q(eoi[5]));
 sky130_fd_sc_hd__dfxtp_2 _27673_ (.CLK(clk),
    .D(_03839_),
    .Q(eoi[6]));
 sky130_fd_sc_hd__dfxtp_2 _27674_ (.CLK(clk),
    .D(_03840_),
    .Q(eoi[7]));
 sky130_fd_sc_hd__dfxtp_2 _27675_ (.CLK(clk),
    .D(_03841_),
    .Q(eoi[8]));
 sky130_fd_sc_hd__dfxtp_2 _27676_ (.CLK(clk),
    .D(_03842_),
    .Q(eoi[9]));
 sky130_fd_sc_hd__dfxtp_2 _27677_ (.CLK(clk),
    .D(_03843_),
    .Q(eoi[10]));
 sky130_fd_sc_hd__dfxtp_2 _27678_ (.CLK(clk),
    .D(_03844_),
    .Q(eoi[11]));
 sky130_fd_sc_hd__dfxtp_2 _27679_ (.CLK(clk),
    .D(_03845_),
    .Q(eoi[12]));
 sky130_fd_sc_hd__dfxtp_2 _27680_ (.CLK(clk),
    .D(_03846_),
    .Q(eoi[13]));
 sky130_fd_sc_hd__dfxtp_2 _27681_ (.CLK(clk),
    .D(_03847_),
    .Q(eoi[14]));
 sky130_fd_sc_hd__dfxtp_2 _27682_ (.CLK(clk),
    .D(_03848_),
    .Q(eoi[15]));
 sky130_fd_sc_hd__dfxtp_2 _27683_ (.CLK(clk),
    .D(_03849_),
    .Q(eoi[16]));
 sky130_fd_sc_hd__dfxtp_2 _27684_ (.CLK(clk),
    .D(_03850_),
    .Q(eoi[17]));
 sky130_fd_sc_hd__dfxtp_2 _27685_ (.CLK(clk),
    .D(_03851_),
    .Q(eoi[18]));
 sky130_fd_sc_hd__dfxtp_2 _27686_ (.CLK(clk),
    .D(_03852_),
    .Q(eoi[19]));
 sky130_fd_sc_hd__dfxtp_2 _27687_ (.CLK(clk),
    .D(_03853_),
    .Q(eoi[20]));
 sky130_fd_sc_hd__dfxtp_2 _27688_ (.CLK(clk),
    .D(_03854_),
    .Q(eoi[21]));
 sky130_fd_sc_hd__dfxtp_2 _27689_ (.CLK(clk),
    .D(_03855_),
    .Q(eoi[22]));
 sky130_fd_sc_hd__dfxtp_2 _27690_ (.CLK(clk),
    .D(_03856_),
    .Q(eoi[23]));
 sky130_fd_sc_hd__dfxtp_2 _27691_ (.CLK(clk),
    .D(_03857_),
    .Q(eoi[24]));
 sky130_fd_sc_hd__dfxtp_2 _27692_ (.CLK(clk),
    .D(_03858_),
    .Q(eoi[25]));
 sky130_fd_sc_hd__dfxtp_2 _27693_ (.CLK(clk),
    .D(_03859_),
    .Q(eoi[26]));
 sky130_fd_sc_hd__dfxtp_2 _27694_ (.CLK(clk),
    .D(_03860_),
    .Q(eoi[27]));
 sky130_fd_sc_hd__dfxtp_2 _27695_ (.CLK(clk),
    .D(_03861_),
    .Q(eoi[28]));
 sky130_fd_sc_hd__dfxtp_2 _27696_ (.CLK(clk),
    .D(_03862_),
    .Q(eoi[29]));
 sky130_fd_sc_hd__dfxtp_2 _27697_ (.CLK(clk),
    .D(_03863_),
    .Q(eoi[30]));
 sky130_fd_sc_hd__dfxtp_2 _27698_ (.CLK(clk),
    .D(_03864_),
    .Q(eoi[31]));
 sky130_fd_sc_hd__dfxtp_2 _27699_ (.CLK(clk),
    .D(_03865_),
    .Q(\count_instr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27700_ (.CLK(clk),
    .D(_03866_),
    .Q(\count_instr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27701_ (.CLK(clk),
    .D(_03867_),
    .Q(\count_instr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27702_ (.CLK(clk),
    .D(_03868_),
    .Q(\count_instr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27703_ (.CLK(clk),
    .D(_03869_),
    .Q(\count_instr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27704_ (.CLK(clk),
    .D(_03870_),
    .Q(\count_instr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27705_ (.CLK(clk),
    .D(_03871_),
    .Q(\count_instr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27706_ (.CLK(clk),
    .D(_03872_),
    .Q(\count_instr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27707_ (.CLK(clk),
    .D(_03873_),
    .Q(\count_instr[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27708_ (.CLK(clk),
    .D(_03874_),
    .Q(\count_instr[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27709_ (.CLK(clk),
    .D(_03875_),
    .Q(\count_instr[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27710_ (.CLK(clk),
    .D(_03876_),
    .Q(\count_instr[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27711_ (.CLK(clk),
    .D(_03877_),
    .Q(\count_instr[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27712_ (.CLK(clk),
    .D(_03878_),
    .Q(\count_instr[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27713_ (.CLK(clk),
    .D(_03879_),
    .Q(\count_instr[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27714_ (.CLK(clk),
    .D(_03880_),
    .Q(\count_instr[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27715_ (.CLK(clk),
    .D(_03881_),
    .Q(\count_instr[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27716_ (.CLK(clk),
    .D(_03882_),
    .Q(\count_instr[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27717_ (.CLK(clk),
    .D(_03883_),
    .Q(\count_instr[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27718_ (.CLK(clk),
    .D(_03884_),
    .Q(\count_instr[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27719_ (.CLK(clk),
    .D(_03885_),
    .Q(\count_instr[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27720_ (.CLK(clk),
    .D(_03886_),
    .Q(\count_instr[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27721_ (.CLK(clk),
    .D(_03887_),
    .Q(\count_instr[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27722_ (.CLK(clk),
    .D(_03888_),
    .Q(\count_instr[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27723_ (.CLK(clk),
    .D(_03889_),
    .Q(\count_instr[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27724_ (.CLK(clk),
    .D(_03890_),
    .Q(\count_instr[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27725_ (.CLK(clk),
    .D(_03891_),
    .Q(\count_instr[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27726_ (.CLK(clk),
    .D(_03892_),
    .Q(\count_instr[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27727_ (.CLK(clk),
    .D(_03893_),
    .Q(\count_instr[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27728_ (.CLK(clk),
    .D(_03894_),
    .Q(\count_instr[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27729_ (.CLK(clk),
    .D(_03895_),
    .Q(\count_instr[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27730_ (.CLK(clk),
    .D(_03896_),
    .Q(\count_instr[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27731_ (.CLK(clk),
    .D(_03897_),
    .Q(\count_instr[32] ));
 sky130_fd_sc_hd__dfxtp_2 _27732_ (.CLK(clk),
    .D(_03898_),
    .Q(\count_instr[33] ));
 sky130_fd_sc_hd__dfxtp_2 _27733_ (.CLK(clk),
    .D(_03899_),
    .Q(\count_instr[34] ));
 sky130_fd_sc_hd__dfxtp_2 _27734_ (.CLK(clk),
    .D(_03900_),
    .Q(\count_instr[35] ));
 sky130_fd_sc_hd__dfxtp_2 _27735_ (.CLK(clk),
    .D(_03901_),
    .Q(\count_instr[36] ));
 sky130_fd_sc_hd__dfxtp_2 _27736_ (.CLK(clk),
    .D(_03902_),
    .Q(\count_instr[37] ));
 sky130_fd_sc_hd__dfxtp_2 _27737_ (.CLK(clk),
    .D(_03903_),
    .Q(\count_instr[38] ));
 sky130_fd_sc_hd__dfxtp_2 _27738_ (.CLK(clk),
    .D(_03904_),
    .Q(\count_instr[39] ));
 sky130_fd_sc_hd__dfxtp_2 _27739_ (.CLK(clk),
    .D(_03905_),
    .Q(\count_instr[40] ));
 sky130_fd_sc_hd__dfxtp_2 _27740_ (.CLK(clk),
    .D(_03906_),
    .Q(\count_instr[41] ));
 sky130_fd_sc_hd__dfxtp_2 _27741_ (.CLK(clk),
    .D(_03907_),
    .Q(\count_instr[42] ));
 sky130_fd_sc_hd__dfxtp_2 _27742_ (.CLK(clk),
    .D(_03908_),
    .Q(\count_instr[43] ));
 sky130_fd_sc_hd__dfxtp_2 _27743_ (.CLK(clk),
    .D(_03909_),
    .Q(\count_instr[44] ));
 sky130_fd_sc_hd__dfxtp_2 _27744_ (.CLK(clk),
    .D(_03910_),
    .Q(\count_instr[45] ));
 sky130_fd_sc_hd__dfxtp_2 _27745_ (.CLK(clk),
    .D(_03911_),
    .Q(\count_instr[46] ));
 sky130_fd_sc_hd__dfxtp_2 _27746_ (.CLK(clk),
    .D(_03912_),
    .Q(\count_instr[47] ));
 sky130_fd_sc_hd__dfxtp_2 _27747_ (.CLK(clk),
    .D(_03913_),
    .Q(\count_instr[48] ));
 sky130_fd_sc_hd__dfxtp_2 _27748_ (.CLK(clk),
    .D(_03914_),
    .Q(\count_instr[49] ));
 sky130_fd_sc_hd__dfxtp_2 _27749_ (.CLK(clk),
    .D(_03915_),
    .Q(\count_instr[50] ));
 sky130_fd_sc_hd__dfxtp_2 _27750_ (.CLK(clk),
    .D(_03916_),
    .Q(\count_instr[51] ));
 sky130_fd_sc_hd__dfxtp_2 _27751_ (.CLK(clk),
    .D(_03917_),
    .Q(\count_instr[52] ));
 sky130_fd_sc_hd__dfxtp_2 _27752_ (.CLK(clk),
    .D(_03918_),
    .Q(\count_instr[53] ));
 sky130_fd_sc_hd__dfxtp_2 _27753_ (.CLK(clk),
    .D(_03919_),
    .Q(\count_instr[54] ));
 sky130_fd_sc_hd__dfxtp_2 _27754_ (.CLK(clk),
    .D(_03920_),
    .Q(\count_instr[55] ));
 sky130_fd_sc_hd__dfxtp_2 _27755_ (.CLK(clk),
    .D(_03921_),
    .Q(\count_instr[56] ));
 sky130_fd_sc_hd__dfxtp_2 _27756_ (.CLK(clk),
    .D(_03922_),
    .Q(\count_instr[57] ));
 sky130_fd_sc_hd__dfxtp_2 _27757_ (.CLK(clk),
    .D(_03923_),
    .Q(\count_instr[58] ));
 sky130_fd_sc_hd__dfxtp_2 _27758_ (.CLK(clk),
    .D(_03924_),
    .Q(\count_instr[59] ));
 sky130_fd_sc_hd__dfxtp_2 _27759_ (.CLK(clk),
    .D(_03925_),
    .Q(\count_instr[60] ));
 sky130_fd_sc_hd__dfxtp_2 _27760_ (.CLK(clk),
    .D(_03926_),
    .Q(\count_instr[61] ));
 sky130_fd_sc_hd__dfxtp_2 _27761_ (.CLK(clk),
    .D(_03927_),
    .Q(\count_instr[62] ));
 sky130_fd_sc_hd__dfxtp_2 _27762_ (.CLK(clk),
    .D(_03928_),
    .Q(\count_instr[63] ));
 sky130_fd_sc_hd__dfxtp_2 _27763_ (.CLK(clk),
    .D(_03929_),
    .Q(\reg_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27764_ (.CLK(clk),
    .D(_03930_),
    .Q(\reg_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27765_ (.CLK(clk),
    .D(_03931_),
    .Q(\reg_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27766_ (.CLK(clk),
    .D(_03932_),
    .Q(\reg_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27767_ (.CLK(clk),
    .D(_03933_),
    .Q(\reg_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27768_ (.CLK(clk),
    .D(_03934_),
    .Q(\reg_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27769_ (.CLK(clk),
    .D(_03935_),
    .Q(\reg_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27770_ (.CLK(clk),
    .D(_03936_),
    .Q(\reg_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27771_ (.CLK(clk),
    .D(_03937_),
    .Q(\reg_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27772_ (.CLK(clk),
    .D(_03938_),
    .Q(\reg_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27773_ (.CLK(clk),
    .D(_03939_),
    .Q(\reg_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27774_ (.CLK(clk),
    .D(_03940_),
    .Q(\reg_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27775_ (.CLK(clk),
    .D(_03941_),
    .Q(\reg_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27776_ (.CLK(clk),
    .D(_03942_),
    .Q(\reg_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27777_ (.CLK(clk),
    .D(_03943_),
    .Q(\reg_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27778_ (.CLK(clk),
    .D(_03944_),
    .Q(\reg_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27779_ (.CLK(clk),
    .D(_03945_),
    .Q(\reg_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27780_ (.CLK(clk),
    .D(_03946_),
    .Q(\reg_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27781_ (.CLK(clk),
    .D(_03947_),
    .Q(\reg_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27782_ (.CLK(clk),
    .D(_03948_),
    .Q(\reg_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27783_ (.CLK(clk),
    .D(_03949_),
    .Q(\reg_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27784_ (.CLK(clk),
    .D(_03950_),
    .Q(\reg_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27785_ (.CLK(clk),
    .D(_03951_),
    .Q(\reg_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27786_ (.CLK(clk),
    .D(_03952_),
    .Q(\reg_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27787_ (.CLK(clk),
    .D(_03953_),
    .Q(\reg_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27788_ (.CLK(clk),
    .D(_03954_),
    .Q(\reg_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27789_ (.CLK(clk),
    .D(_03955_),
    .Q(\reg_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27790_ (.CLK(clk),
    .D(_03956_),
    .Q(\reg_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27791_ (.CLK(clk),
    .D(_03957_),
    .Q(\reg_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27792_ (.CLK(clk),
    .D(_03958_),
    .Q(\reg_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27793_ (.CLK(clk),
    .D(_03959_),
    .Q(\reg_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27794_ (.CLK(clk),
    .D(_03960_),
    .Q(\reg_next_pc[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27795_ (.CLK(clk),
    .D(_03961_),
    .Q(\reg_next_pc[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27796_ (.CLK(clk),
    .D(_03962_),
    .Q(\reg_next_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27797_ (.CLK(clk),
    .D(_03963_),
    .Q(\reg_next_pc[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27798_ (.CLK(clk),
    .D(_03964_),
    .Q(\reg_next_pc[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27799_ (.CLK(clk),
    .D(_03965_),
    .Q(\reg_next_pc[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27800_ (.CLK(clk),
    .D(_03966_),
    .Q(\reg_next_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27801_ (.CLK(clk),
    .D(_03967_),
    .Q(\reg_next_pc[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27802_ (.CLK(clk),
    .D(_03968_),
    .Q(\reg_next_pc[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27803_ (.CLK(clk),
    .D(_03969_),
    .Q(\reg_next_pc[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27804_ (.CLK(clk),
    .D(_03970_),
    .Q(\reg_next_pc[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27805_ (.CLK(clk),
    .D(_03971_),
    .Q(\reg_next_pc[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27806_ (.CLK(clk),
    .D(_03972_),
    .Q(\reg_next_pc[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27807_ (.CLK(clk),
    .D(_03973_),
    .Q(\reg_next_pc[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27808_ (.CLK(clk),
    .D(_03974_),
    .Q(\reg_next_pc[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27809_ (.CLK(clk),
    .D(_03975_),
    .Q(\reg_next_pc[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27810_ (.CLK(clk),
    .D(_03976_),
    .Q(\reg_next_pc[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27811_ (.CLK(clk),
    .D(_03977_),
    .Q(\reg_next_pc[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27812_ (.CLK(clk),
    .D(_03978_),
    .Q(\reg_next_pc[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27813_ (.CLK(clk),
    .D(_03979_),
    .Q(\reg_next_pc[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27814_ (.CLK(clk),
    .D(_03980_),
    .Q(\reg_next_pc[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27815_ (.CLK(clk),
    .D(_03981_),
    .Q(\reg_next_pc[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27816_ (.CLK(clk),
    .D(_03982_),
    .Q(\reg_next_pc[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27817_ (.CLK(clk),
    .D(_03983_),
    .Q(\reg_next_pc[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27818_ (.CLK(clk),
    .D(_03984_),
    .Q(\reg_next_pc[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27819_ (.CLK(clk),
    .D(_03985_),
    .Q(\reg_next_pc[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27820_ (.CLK(clk),
    .D(_03986_),
    .Q(\reg_next_pc[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27821_ (.CLK(clk),
    .D(_03987_),
    .Q(\reg_next_pc[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27822_ (.CLK(clk),
    .D(_03988_),
    .Q(\reg_next_pc[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27823_ (.CLK(clk),
    .D(_03989_),
    .Q(\reg_next_pc[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27824_ (.CLK(clk),
    .D(_03990_),
    .Q(\reg_next_pc[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27825_ (.CLK(clk),
    .D(_03991_),
    .Q(mem_do_rdata));
 sky130_fd_sc_hd__dfxtp_2 _27826_ (.CLK(clk),
    .D(_03992_),
    .Q(mem_do_wdata));
 sky130_fd_sc_hd__dfxtp_2 _27827_ (.CLK(clk),
    .D(_03993_),
    .Q(\pcpi_timeout_counter[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27828_ (.CLK(clk),
    .D(_03994_),
    .Q(\pcpi_timeout_counter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27829_ (.CLK(clk),
    .D(_03995_),
    .Q(\pcpi_timeout_counter[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27830_ (.CLK(clk),
    .D(_03996_),
    .Q(\pcpi_timeout_counter[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27831_ (.CLK(clk),
    .D(_03997_),
    .Q(instr_beq));
 sky130_fd_sc_hd__dfxtp_2 _27832_ (.CLK(clk),
    .D(_03998_),
    .Q(instr_bne));
 sky130_fd_sc_hd__dfxtp_2 _27833_ (.CLK(clk),
    .D(_03999_),
    .Q(instr_blt));
 sky130_fd_sc_hd__dfxtp_2 _27834_ (.CLK(clk),
    .D(_04000_),
    .Q(instr_bge));
 sky130_fd_sc_hd__dfxtp_2 _27835_ (.CLK(clk),
    .D(_04001_),
    .Q(instr_bltu));
 sky130_fd_sc_hd__dfxtp_2 _27836_ (.CLK(clk),
    .D(_04002_),
    .Q(instr_bgeu));
 sky130_fd_sc_hd__dfxtp_2 _27837_ (.CLK(clk),
    .D(_04003_),
    .Q(instr_addi));
 sky130_fd_sc_hd__dfxtp_2 _27838_ (.CLK(clk),
    .D(_04004_),
    .Q(instr_slti));
 sky130_fd_sc_hd__dfxtp_2 _27839_ (.CLK(clk),
    .D(_04005_),
    .Q(instr_sltiu));
 sky130_fd_sc_hd__dfxtp_2 _27840_ (.CLK(clk),
    .D(_04006_),
    .Q(instr_xori));
 sky130_fd_sc_hd__dfxtp_2 _27841_ (.CLK(clk),
    .D(_04007_),
    .Q(instr_ori));
 sky130_fd_sc_hd__dfxtp_2 _27842_ (.CLK(clk),
    .D(_04008_),
    .Q(instr_andi));
 sky130_fd_sc_hd__dfxtp_2 _27843_ (.CLK(clk),
    .D(_04009_),
    .Q(instr_add));
 sky130_fd_sc_hd__dfxtp_2 _27844_ (.CLK(clk),
    .D(_04010_),
    .Q(instr_sub));
 sky130_fd_sc_hd__dfxtp_2 _27845_ (.CLK(clk),
    .D(_04011_),
    .Q(instr_sll));
 sky130_fd_sc_hd__dfxtp_2 _27846_ (.CLK(clk),
    .D(_04012_),
    .Q(instr_slt));
 sky130_fd_sc_hd__dfxtp_2 _27847_ (.CLK(clk),
    .D(_04013_),
    .Q(instr_sltu));
 sky130_fd_sc_hd__dfxtp_2 _27848_ (.CLK(clk),
    .D(_04014_),
    .Q(instr_xor));
 sky130_fd_sc_hd__dfxtp_2 _27849_ (.CLK(clk),
    .D(_04015_),
    .Q(instr_srl));
 sky130_fd_sc_hd__dfxtp_2 _27850_ (.CLK(clk),
    .D(_04016_),
    .Q(instr_sra));
 sky130_fd_sc_hd__dfxtp_2 _27851_ (.CLK(clk),
    .D(_04017_),
    .Q(instr_or));
 sky130_fd_sc_hd__dfxtp_2 _27852_ (.CLK(clk),
    .D(_04018_),
    .Q(instr_and));
 sky130_fd_sc_hd__dfxtp_2 _27853_ (.CLK(clk),
    .D(_04019_),
    .Q(\decoded_rs1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27854_ (.CLK(clk),
    .D(_04020_),
    .Q(\decoded_rs1[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27855_ (.CLK(clk),
    .D(_04021_),
    .Q(\decoded_rs1[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27856_ (.CLK(clk),
    .D(_04022_),
    .Q(\decoded_rs1[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27857_ (.CLK(clk),
    .D(_04023_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu));
 sky130_fd_sc_hd__dfxtp_2 _27858_ (.CLK(clk),
    .D(_04024_),
    .Q(mem_instr));
 sky130_fd_sc_hd__dfxtp_2 _27859_ (.CLK(clk),
    .D(_04025_),
    .Q(\irq_mask[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27860_ (.CLK(clk),
    .D(_04026_),
    .Q(\irq_mask[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27861_ (.CLK(clk),
    .D(_04027_),
    .Q(\irq_mask[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27862_ (.CLK(clk),
    .D(_04028_),
    .Q(\irq_mask[3] ));
 sky130_fd_sc_hd__dfxtp_2 _27863_ (.CLK(clk),
    .D(_04029_),
    .Q(\irq_mask[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27864_ (.CLK(clk),
    .D(_04030_),
    .Q(\irq_mask[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27865_ (.CLK(clk),
    .D(_04031_),
    .Q(\irq_mask[6] ));
 sky130_fd_sc_hd__dfxtp_2 _27866_ (.CLK(clk),
    .D(_04032_),
    .Q(\irq_mask[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27867_ (.CLK(clk),
    .D(_04033_),
    .Q(\irq_mask[8] ));
 sky130_fd_sc_hd__dfxtp_2 _27868_ (.CLK(clk),
    .D(_04034_),
    .Q(\irq_mask[9] ));
 sky130_fd_sc_hd__dfxtp_2 _27869_ (.CLK(clk),
    .D(_04035_),
    .Q(\irq_mask[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27870_ (.CLK(clk),
    .D(_04036_),
    .Q(\irq_mask[11] ));
 sky130_fd_sc_hd__dfxtp_2 _27871_ (.CLK(clk),
    .D(_04037_),
    .Q(\irq_mask[12] ));
 sky130_fd_sc_hd__dfxtp_2 _27872_ (.CLK(clk),
    .D(_04038_),
    .Q(\irq_mask[13] ));
 sky130_fd_sc_hd__dfxtp_2 _27873_ (.CLK(clk),
    .D(_04039_),
    .Q(\irq_mask[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27874_ (.CLK(clk),
    .D(_04040_),
    .Q(\irq_mask[15] ));
 sky130_fd_sc_hd__dfxtp_2 _27875_ (.CLK(clk),
    .D(_04041_),
    .Q(\irq_mask[16] ));
 sky130_fd_sc_hd__dfxtp_2 _27876_ (.CLK(clk),
    .D(_04042_),
    .Q(\irq_mask[17] ));
 sky130_fd_sc_hd__dfxtp_2 _27877_ (.CLK(clk),
    .D(_04043_),
    .Q(\irq_mask[18] ));
 sky130_fd_sc_hd__dfxtp_2 _27878_ (.CLK(clk),
    .D(_04044_),
    .Q(\irq_mask[19] ));
 sky130_fd_sc_hd__dfxtp_2 _27879_ (.CLK(clk),
    .D(_04045_),
    .Q(\irq_mask[20] ));
 sky130_fd_sc_hd__dfxtp_2 _27880_ (.CLK(clk),
    .D(_04046_),
    .Q(\irq_mask[21] ));
 sky130_fd_sc_hd__dfxtp_2 _27881_ (.CLK(clk),
    .D(_04047_),
    .Q(\irq_mask[22] ));
 sky130_fd_sc_hd__dfxtp_2 _27882_ (.CLK(clk),
    .D(_04048_),
    .Q(\irq_mask[23] ));
 sky130_fd_sc_hd__dfxtp_2 _27883_ (.CLK(clk),
    .D(_04049_),
    .Q(\irq_mask[24] ));
 sky130_fd_sc_hd__dfxtp_2 _27884_ (.CLK(clk),
    .D(_04050_),
    .Q(\irq_mask[25] ));
 sky130_fd_sc_hd__dfxtp_2 _27885_ (.CLK(clk),
    .D(_04051_),
    .Q(\irq_mask[26] ));
 sky130_fd_sc_hd__dfxtp_2 _27886_ (.CLK(clk),
    .D(_04052_),
    .Q(\irq_mask[27] ));
 sky130_fd_sc_hd__dfxtp_2 _27887_ (.CLK(clk),
    .D(_04053_),
    .Q(\irq_mask[28] ));
 sky130_fd_sc_hd__dfxtp_2 _27888_ (.CLK(clk),
    .D(_04054_),
    .Q(\irq_mask[29] ));
 sky130_fd_sc_hd__dfxtp_2 _27889_ (.CLK(clk),
    .D(_04055_),
    .Q(\irq_mask[30] ));
 sky130_fd_sc_hd__dfxtp_2 _27890_ (.CLK(clk),
    .D(_04056_),
    .Q(\irq_mask[31] ));
 sky130_fd_sc_hd__dfxtp_2 _27891_ (.CLK(clk),
    .D(_04057_),
    .Q(mem_do_prefetch));
 sky130_fd_sc_hd__dfxtp_2 _27892_ (.CLK(clk),
    .D(_04058_),
    .Q(mem_do_rinst));
 sky130_fd_sc_hd__dfxtp_2 _27893_ (.CLK(clk),
    .D(_04059_),
    .Q(\irq_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27894_ (.CLK(clk),
    .D(_04060_),
    .Q(\irq_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27895_ (.CLK(clk),
    .D(_04061_),
    .Q(latched_store));
 sky130_fd_sc_hd__dfxtp_2 _27896_ (.CLK(clk),
    .D(_04062_),
    .Q(latched_stalu));
 sky130_fd_sc_hd__dfxtp_2 _27897_ (.CLK(clk),
    .D(_04063_),
    .Q(\pcpi_mul.rs2[32] ));
 sky130_fd_sc_hd__dfxtp_2 _27898_ (.CLK(clk),
    .D(_04064_),
    .Q(\pcpi_mul.rs1[32] ));
 sky130_fd_sc_hd__dfxtp_2 _27899_ (.CLK(clk),
    .D(_04065_),
    .Q(irq_delay));
 sky130_fd_sc_hd__dfxtp_2 _27900_ (.CLK(clk),
    .D(_04066_),
    .Q(\decoded_rs1[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27901_ (.CLK(clk),
    .D(_04067_),
    .Q(\mem_state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27902_ (.CLK(clk),
    .D(_04068_),
    .Q(\mem_state[1] ));
 sky130_fd_sc_hd__dfxtp_2 _27903_ (.CLK(clk),
    .D(_04069_),
    .Q(latched_branch));
 sky130_fd_sc_hd__dfxtp_2 _27904_ (.CLK(clk),
    .D(_04070_),
    .Q(latched_is_lh));
 sky130_fd_sc_hd__dfxtp_2 _27905_ (.CLK(clk),
    .D(_04071_),
    .Q(latched_is_lb));
 sky130_fd_sc_hd__dfxtp_2 _27906_ (.CLK(clk),
    .D(_04072_),
    .Q(irq_active));
endmodule
